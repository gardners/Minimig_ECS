library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

--
entity audio_data is
  port (ClkA : in std_logic;
        addressa : in integer range 0 to 65535;
        doa : out std_logic_vector(7 downto 0)
        );
end audio_data;

architecture Behavioral of audio_data is

  type ram_t is array (0 to 65535) of std_logic_vector(7 downto 0);
  shared variable ram : ram_t := (
          0 => x"52", -- $00000
          1 => x"49", -- $00001
          2 => x"46", -- $00002
          3 => x"46", -- $00003
          4 => x"46", -- $00004
          5 => x"ac", -- $00005
          6 => x"00", -- $00006
          7 => x"00", -- $00007
          8 => x"57", -- $00008
          9 => x"41", -- $00009
          10 => x"56", -- $0000a
          11 => x"45", -- $0000b
          12 => x"66", -- $0000c
          13 => x"6d", -- $0000d
          14 => x"74", -- $0000e
          15 => x"20", -- $0000f
          16 => x"10", -- $00010
          17 => x"00", -- $00011
          18 => x"00", -- $00012
          19 => x"00", -- $00013
          20 => x"01", -- $00014
          21 => x"00", -- $00015
          22 => x"01", -- $00016
          23 => x"00", -- $00017
          24 => x"40", -- $00018
          25 => x"1f", -- $00019
          26 => x"00", -- $0001a
          27 => x"00", -- $0001b
          28 => x"40", -- $0001c
          29 => x"1f", -- $0001d
          30 => x"00", -- $0001e
          31 => x"00", -- $0001f
          32 => x"01", -- $00020
          33 => x"00", -- $00021
          34 => x"08", -- $00022
          35 => x"00", -- $00023
          36 => x"4c", -- $00024
          37 => x"49", -- $00025
          38 => x"53", -- $00026
          39 => x"54", -- $00027
          40 => x"1a", -- $00028
          41 => x"00", -- $00029
          42 => x"00", -- $0002a
          43 => x"00", -- $0002b
          44 => x"49", -- $0002c
          45 => x"4e", -- $0002d
          46 => x"46", -- $0002e
          47 => x"4f", -- $0002f
          48 => x"49", -- $00030
          49 => x"53", -- $00031
          50 => x"46", -- $00032
          51 => x"54", -- $00033
          52 => x"0e", -- $00034
          53 => x"00", -- $00035
          54 => x"00", -- $00036
          55 => x"00", -- $00037
          56 => x"4c", -- $00038
          57 => x"61", -- $00039
          58 => x"76", -- $0003a
          59 => x"66", -- $0003b
          60 => x"35", -- $0003c
          61 => x"37", -- $0003d
          62 => x"2e", -- $0003e
          63 => x"38", -- $0003f
          64 => x"33", -- $00040
          65 => x"2e", -- $00041
          66 => x"31", -- $00042
          67 => x"30", -- $00043
          68 => x"30", -- $00044
          69 => x"00", -- $00045
          70 => x"64", -- $00046
          71 => x"61", -- $00047
          72 => x"74", -- $00048
          73 => x"61", -- $00049
          74 => x"00", -- $0004a
          75 => x"ac", -- $0004b
          76 => x"00", -- $0004c
          77 => x"00", -- $0004d
          78 => x"80", -- $0004e
          79 => x"80", -- $0004f
          80 => x"80", -- $00050
          81 => x"80", -- $00051
          82 => x"80", -- $00052
          83 => x"80", -- $00053
          84 => x"80", -- $00054
          85 => x"80", -- $00055
          86 => x"80", -- $00056
          87 => x"80", -- $00057
          88 => x"80", -- $00058
          89 => x"80", -- $00059
          90 => x"80", -- $0005a
          91 => x"80", -- $0005b
          92 => x"80", -- $0005c
          93 => x"80", -- $0005d
          94 => x"80", -- $0005e
          95 => x"80", -- $0005f
          96 => x"80", -- $00060
          97 => x"80", -- $00061
          98 => x"80", -- $00062
          99 => x"80", -- $00063
          100 => x"80", -- $00064
          101 => x"80", -- $00065
          102 => x"80", -- $00066
          103 => x"80", -- $00067
          104 => x"80", -- $00068
          105 => x"80", -- $00069
          106 => x"80", -- $0006a
          107 => x"80", -- $0006b
          108 => x"80", -- $0006c
          109 => x"80", -- $0006d
          110 => x"80", -- $0006e
          111 => x"80", -- $0006f
          112 => x"80", -- $00070
          113 => x"80", -- $00071
          114 => x"80", -- $00072
          115 => x"80", -- $00073
          116 => x"80", -- $00074
          117 => x"80", -- $00075
          118 => x"80", -- $00076
          119 => x"7f", -- $00077
          120 => x"7f", -- $00078
          121 => x"7f", -- $00079
          122 => x"7f", -- $0007a
          123 => x"7f", -- $0007b
          124 => x"80", -- $0007c
          125 => x"80", -- $0007d
          126 => x"80", -- $0007e
          127 => x"80", -- $0007f
          128 => x"80", -- $00080
          129 => x"80", -- $00081
          130 => x"80", -- $00082
          131 => x"80", -- $00083
          132 => x"80", -- $00084
          133 => x"80", -- $00085
          134 => x"7f", -- $00086
          135 => x"7f", -- $00087
          136 => x"7f", -- $00088
          137 => x"7f", -- $00089
          138 => x"7f", -- $0008a
          139 => x"7f", -- $0008b
          140 => x"7f", -- $0008c
          141 => x"7f", -- $0008d
          142 => x"7f", -- $0008e
          143 => x"7f", -- $0008f
          144 => x"7f", -- $00090
          145 => x"7f", -- $00091
          146 => x"7f", -- $00092
          147 => x"7f", -- $00093
          148 => x"7f", -- $00094
          149 => x"7f", -- $00095
          150 => x"7f", -- $00096
          151 => x"7f", -- $00097
          152 => x"7f", -- $00098
          153 => x"7e", -- $00099
          154 => x"7e", -- $0009a
          155 => x"7e", -- $0009b
          156 => x"7e", -- $0009c
          157 => x"7e", -- $0009d
          158 => x"7e", -- $0009e
          159 => x"7e", -- $0009f
          160 => x"7e", -- $000a0
          161 => x"7e", -- $000a1
          162 => x"7d", -- $000a2
          163 => x"7d", -- $000a3
          164 => x"7d", -- $000a4
          165 => x"7d", -- $000a5
          166 => x"7d", -- $000a6
          167 => x"7d", -- $000a7
          168 => x"7d", -- $000a8
          169 => x"7d", -- $000a9
          170 => x"7d", -- $000aa
          171 => x"7d", -- $000ab
          172 => x"7d", -- $000ac
          173 => x"7d", -- $000ad
          174 => x"7d", -- $000ae
          175 => x"7d", -- $000af
          176 => x"7d", -- $000b0
          177 => x"7d", -- $000b1
          178 => x"7d", -- $000b2
          179 => x"7d", -- $000b3
          180 => x"7d", -- $000b4
          181 => x"7d", -- $000b5
          182 => x"7d", -- $000b6
          183 => x"7d", -- $000b7
          184 => x"7d", -- $000b8
          185 => x"7d", -- $000b9
          186 => x"7d", -- $000ba
          187 => x"7c", -- $000bb
          188 => x"7d", -- $000bc
          189 => x"7d", -- $000bd
          190 => x"7d", -- $000be
          191 => x"7d", -- $000bf
          192 => x"7d", -- $000c0
          193 => x"7d", -- $000c1
          194 => x"7c", -- $000c2
          195 => x"7c", -- $000c3
          196 => x"7c", -- $000c4
          197 => x"7d", -- $000c5
          198 => x"7d", -- $000c6
          199 => x"7d", -- $000c7
          200 => x"7c", -- $000c8
          201 => x"7c", -- $000c9
          202 => x"7c", -- $000ca
          203 => x"7d", -- $000cb
          204 => x"7c", -- $000cc
          205 => x"7d", -- $000cd
          206 => x"7d", -- $000ce
          207 => x"7d", -- $000cf
          208 => x"7d", -- $000d0
          209 => x"7d", -- $000d1
          210 => x"7d", -- $000d2
          211 => x"7d", -- $000d3
          212 => x"7d", -- $000d4
          213 => x"7d", -- $000d5
          214 => x"7d", -- $000d6
          215 => x"7d", -- $000d7
          216 => x"7d", -- $000d8
          217 => x"7d", -- $000d9
          218 => x"7d", -- $000da
          219 => x"7d", -- $000db
          220 => x"7d", -- $000dc
          221 => x"7d", -- $000dd
          222 => x"7d", -- $000de
          223 => x"7d", -- $000df
          224 => x"7d", -- $000e0
          225 => x"7d", -- $000e1
          226 => x"7d", -- $000e2
          227 => x"7d", -- $000e3
          228 => x"7d", -- $000e4
          229 => x"7d", -- $000e5
          230 => x"7d", -- $000e6
          231 => x"7d", -- $000e7
          232 => x"7d", -- $000e8
          233 => x"7d", -- $000e9
          234 => x"7d", -- $000ea
          235 => x"7d", -- $000eb
          236 => x"7d", -- $000ec
          237 => x"7d", -- $000ed
          238 => x"7d", -- $000ee
          239 => x"7d", -- $000ef
          240 => x"7d", -- $000f0
          241 => x"7d", -- $000f1
          242 => x"7d", -- $000f2
          243 => x"7d", -- $000f3
          244 => x"7d", -- $000f4
          245 => x"7d", -- $000f5
          246 => x"7d", -- $000f6
          247 => x"7d", -- $000f7
          248 => x"7d", -- $000f8
          249 => x"7d", -- $000f9
          250 => x"7d", -- $000fa
          251 => x"7c", -- $000fb
          252 => x"7c", -- $000fc
          253 => x"7c", -- $000fd
          254 => x"7c", -- $000fe
          255 => x"7c", -- $000ff
          256 => x"7c", -- $00100
          257 => x"7c", -- $00101
          258 => x"7c", -- $00102
          259 => x"7c", -- $00103
          260 => x"7c", -- $00104
          261 => x"7c", -- $00105
          262 => x"7c", -- $00106
          263 => x"7c", -- $00107
          264 => x"7c", -- $00108
          265 => x"7c", -- $00109
          266 => x"7c", -- $0010a
          267 => x"7c", -- $0010b
          268 => x"7c", -- $0010c
          269 => x"7c", -- $0010d
          270 => x"7c", -- $0010e
          271 => x"7c", -- $0010f
          272 => x"7b", -- $00110
          273 => x"7c", -- $00111
          274 => x"7b", -- $00112
          275 => x"7c", -- $00113
          276 => x"7c", -- $00114
          277 => x"7c", -- $00115
          278 => x"7c", -- $00116
          279 => x"7b", -- $00117
          280 => x"7b", -- $00118
          281 => x"7b", -- $00119
          282 => x"7b", -- $0011a
          283 => x"7b", -- $0011b
          284 => x"7c", -- $0011c
          285 => x"7b", -- $0011d
          286 => x"7b", -- $0011e
          287 => x"7b", -- $0011f
          288 => x"7b", -- $00120
          289 => x"7b", -- $00121
          290 => x"7b", -- $00122
          291 => x"7b", -- $00123
          292 => x"7b", -- $00124
          293 => x"7b", -- $00125
          294 => x"7b", -- $00126
          295 => x"7b", -- $00127
          296 => x"7b", -- $00128
          297 => x"7b", -- $00129
          298 => x"7b", -- $0012a
          299 => x"7b", -- $0012b
          300 => x"7b", -- $0012c
          301 => x"7b", -- $0012d
          302 => x"7b", -- $0012e
          303 => x"7b", -- $0012f
          304 => x"7b", -- $00130
          305 => x"7b", -- $00131
          306 => x"7b", -- $00132
          307 => x"7b", -- $00133
          308 => x"7b", -- $00134
          309 => x"7b", -- $00135
          310 => x"7b", -- $00136
          311 => x"7b", -- $00137
          312 => x"7b", -- $00138
          313 => x"7b", -- $00139
          314 => x"7b", -- $0013a
          315 => x"7b", -- $0013b
          316 => x"7b", -- $0013c
          317 => x"7b", -- $0013d
          318 => x"7b", -- $0013e
          319 => x"7b", -- $0013f
          320 => x"7c", -- $00140
          321 => x"7b", -- $00141
          322 => x"7b", -- $00142
          323 => x"7b", -- $00143
          324 => x"7b", -- $00144
          325 => x"7c", -- $00145
          326 => x"7c", -- $00146
          327 => x"7c", -- $00147
          328 => x"7c", -- $00148
          329 => x"7c", -- $00149
          330 => x"7c", -- $0014a
          331 => x"7c", -- $0014b
          332 => x"7c", -- $0014c
          333 => x"7b", -- $0014d
          334 => x"7b", -- $0014e
          335 => x"7c", -- $0014f
          336 => x"7c", -- $00150
          337 => x"7c", -- $00151
          338 => x"7c", -- $00152
          339 => x"7c", -- $00153
          340 => x"7b", -- $00154
          341 => x"7b", -- $00155
          342 => x"7c", -- $00156
          343 => x"7c", -- $00157
          344 => x"7c", -- $00158
          345 => x"7c", -- $00159
          346 => x"7c", -- $0015a
          347 => x"7b", -- $0015b
          348 => x"7b", -- $0015c
          349 => x"7c", -- $0015d
          350 => x"7c", -- $0015e
          351 => x"7c", -- $0015f
          352 => x"7c", -- $00160
          353 => x"7c", -- $00161
          354 => x"7c", -- $00162
          355 => x"7c", -- $00163
          356 => x"7c", -- $00164
          357 => x"7c", -- $00165
          358 => x"7c", -- $00166
          359 => x"7c", -- $00167
          360 => x"7c", -- $00168
          361 => x"7c", -- $00169
          362 => x"7c", -- $0016a
          363 => x"7c", -- $0016b
          364 => x"7c", -- $0016c
          365 => x"7c", -- $0016d
          366 => x"7c", -- $0016e
          367 => x"7c", -- $0016f
          368 => x"7c", -- $00170
          369 => x"7c", -- $00171
          370 => x"7c", -- $00172
          371 => x"7c", -- $00173
          372 => x"7c", -- $00174
          373 => x"7c", -- $00175
          374 => x"7c", -- $00176
          375 => x"7c", -- $00177
          376 => x"7c", -- $00178
          377 => x"7d", -- $00179
          378 => x"7d", -- $0017a
          379 => x"7c", -- $0017b
          380 => x"7c", -- $0017c
          381 => x"7c", -- $0017d
          382 => x"7c", -- $0017e
          383 => x"7c", -- $0017f
          384 => x"7c", -- $00180
          385 => x"7d", -- $00181
          386 => x"7d", -- $00182
          387 => x"7d", -- $00183
          388 => x"7d", -- $00184
          389 => x"7d", -- $00185
          390 => x"7d", -- $00186
          391 => x"7d", -- $00187
          392 => x"7d", -- $00188
          393 => x"7d", -- $00189
          394 => x"7d", -- $0018a
          395 => x"7d", -- $0018b
          396 => x"7d", -- $0018c
          397 => x"7d", -- $0018d
          398 => x"7d", -- $0018e
          399 => x"7d", -- $0018f
          400 => x"7d", -- $00190
          401 => x"7d", -- $00191
          402 => x"7e", -- $00192
          403 => x"7e", -- $00193
          404 => x"7d", -- $00194
          405 => x"7d", -- $00195
          406 => x"7d", -- $00196
          407 => x"7e", -- $00197
          408 => x"7e", -- $00198
          409 => x"7e", -- $00199
          410 => x"7e", -- $0019a
          411 => x"7e", -- $0019b
          412 => x"7e", -- $0019c
          413 => x"7e", -- $0019d
          414 => x"7e", -- $0019e
          415 => x"7e", -- $0019f
          416 => x"7e", -- $001a0
          417 => x"7e", -- $001a1
          418 => x"7e", -- $001a2
          419 => x"7e", -- $001a3
          420 => x"7e", -- $001a4
          421 => x"7e", -- $001a5
          422 => x"7e", -- $001a6
          423 => x"7e", -- $001a7
          424 => x"7e", -- $001a8
          425 => x"7f", -- $001a9
          426 => x"7f", -- $001aa
          427 => x"7f", -- $001ab
          428 => x"7f", -- $001ac
          429 => x"7f", -- $001ad
          430 => x"7f", -- $001ae
          431 => x"7e", -- $001af
          432 => x"7f", -- $001b0
          433 => x"7f", -- $001b1
          434 => x"7f", -- $001b2
          435 => x"7f", -- $001b3
          436 => x"7f", -- $001b4
          437 => x"7f", -- $001b5
          438 => x"7f", -- $001b6
          439 => x"7f", -- $001b7
          440 => x"7f", -- $001b8
          441 => x"7f", -- $001b9
          442 => x"7f", -- $001ba
          443 => x"7f", -- $001bb
          444 => x"7f", -- $001bc
          445 => x"7f", -- $001bd
          446 => x"80", -- $001be
          447 => x"80", -- $001bf
          448 => x"80", -- $001c0
          449 => x"80", -- $001c1
          450 => x"80", -- $001c2
          451 => x"80", -- $001c3
          452 => x"80", -- $001c4
          453 => x"80", -- $001c5
          454 => x"80", -- $001c6
          455 => x"80", -- $001c7
          456 => x"80", -- $001c8
          457 => x"80", -- $001c9
          458 => x"80", -- $001ca
          459 => x"80", -- $001cb
          460 => x"80", -- $001cc
          461 => x"80", -- $001cd
          462 => x"80", -- $001ce
          463 => x"80", -- $001cf
          464 => x"80", -- $001d0
          465 => x"80", -- $001d1
          466 => x"80", -- $001d2
          467 => x"80", -- $001d3
          468 => x"80", -- $001d4
          469 => x"80", -- $001d5
          470 => x"81", -- $001d6
          471 => x"81", -- $001d7
          472 => x"81", -- $001d8
          473 => x"81", -- $001d9
          474 => x"81", -- $001da
          475 => x"81", -- $001db
          476 => x"81", -- $001dc
          477 => x"81", -- $001dd
          478 => x"81", -- $001de
          479 => x"81", -- $001df
          480 => x"81", -- $001e0
          481 => x"81", -- $001e1
          482 => x"81", -- $001e2
          483 => x"81", -- $001e3
          484 => x"81", -- $001e4
          485 => x"81", -- $001e5
          486 => x"81", -- $001e6
          487 => x"81", -- $001e7
          488 => x"81", -- $001e8
          489 => x"81", -- $001e9
          490 => x"81", -- $001ea
          491 => x"81", -- $001eb
          492 => x"81", -- $001ec
          493 => x"81", -- $001ed
          494 => x"81", -- $001ee
          495 => x"82", -- $001ef
          496 => x"82", -- $001f0
          497 => x"82", -- $001f1
          498 => x"82", -- $001f2
          499 => x"81", -- $001f3
          500 => x"81", -- $001f4
          501 => x"82", -- $001f5
          502 => x"82", -- $001f6
          503 => x"82", -- $001f7
          504 => x"82", -- $001f8
          505 => x"82", -- $001f9
          506 => x"82", -- $001fa
          507 => x"82", -- $001fb
          508 => x"82", -- $001fc
          509 => x"82", -- $001fd
          510 => x"82", -- $001fe
          511 => x"82", -- $001ff
          512 => x"82", -- $00200
          513 => x"82", -- $00201
          514 => x"82", -- $00202
          515 => x"82", -- $00203
          516 => x"82", -- $00204
          517 => x"82", -- $00205
          518 => x"82", -- $00206
          519 => x"82", -- $00207
          520 => x"82", -- $00208
          521 => x"83", -- $00209
          522 => x"83", -- $0020a
          523 => x"82", -- $0020b
          524 => x"82", -- $0020c
          525 => x"82", -- $0020d
          526 => x"82", -- $0020e
          527 => x"82", -- $0020f
          528 => x"82", -- $00210
          529 => x"82", -- $00211
          530 => x"82", -- $00212
          531 => x"82", -- $00213
          532 => x"82", -- $00214
          533 => x"82", -- $00215
          534 => x"82", -- $00216
          535 => x"82", -- $00217
          536 => x"82", -- $00218
          537 => x"82", -- $00219
          538 => x"82", -- $0021a
          539 => x"82", -- $0021b
          540 => x"82", -- $0021c
          541 => x"82", -- $0021d
          542 => x"82", -- $0021e
          543 => x"82", -- $0021f
          544 => x"83", -- $00220
          545 => x"83", -- $00221
          546 => x"83", -- $00222
          547 => x"83", -- $00223
          548 => x"82", -- $00224
          549 => x"82", -- $00225
          550 => x"82", -- $00226
          551 => x"82", -- $00227
          552 => x"83", -- $00228
          553 => x"83", -- $00229
          554 => x"83", -- $0022a
          555 => x"82", -- $0022b
          556 => x"83", -- $0022c
          557 => x"83", -- $0022d
          558 => x"83", -- $0022e
          559 => x"83", -- $0022f
          560 => x"83", -- $00230
          561 => x"83", -- $00231
          562 => x"83", -- $00232
          563 => x"83", -- $00233
          564 => x"83", -- $00234
          565 => x"83", -- $00235
          566 => x"83", -- $00236
          567 => x"83", -- $00237
          568 => x"83", -- $00238
          569 => x"83", -- $00239
          570 => x"83", -- $0023a
          571 => x"83", -- $0023b
          572 => x"83", -- $0023c
          573 => x"83", -- $0023d
          574 => x"83", -- $0023e
          575 => x"83", -- $0023f
          576 => x"83", -- $00240
          577 => x"83", -- $00241
          578 => x"83", -- $00242
          579 => x"83", -- $00243
          580 => x"83", -- $00244
          581 => x"83", -- $00245
          582 => x"83", -- $00246
          583 => x"83", -- $00247
          584 => x"83", -- $00248
          585 => x"83", -- $00249
          586 => x"83", -- $0024a
          587 => x"83", -- $0024b
          588 => x"83", -- $0024c
          589 => x"83", -- $0024d
          590 => x"83", -- $0024e
          591 => x"83", -- $0024f
          592 => x"83", -- $00250
          593 => x"84", -- $00251
          594 => x"84", -- $00252
          595 => x"84", -- $00253
          596 => x"84", -- $00254
          597 => x"84", -- $00255
          598 => x"84", -- $00256
          599 => x"83", -- $00257
          600 => x"84", -- $00258
          601 => x"84", -- $00259
          602 => x"84", -- $0025a
          603 => x"84", -- $0025b
          604 => x"84", -- $0025c
          605 => x"84", -- $0025d
          606 => x"84", -- $0025e
          607 => x"84", -- $0025f
          608 => x"84", -- $00260
          609 => x"84", -- $00261
          610 => x"84", -- $00262
          611 => x"84", -- $00263
          612 => x"84", -- $00264
          613 => x"84", -- $00265
          614 => x"84", -- $00266
          615 => x"84", -- $00267
          616 => x"84", -- $00268
          617 => x"84", -- $00269
          618 => x"85", -- $0026a
          619 => x"85", -- $0026b
          620 => x"85", -- $0026c
          621 => x"85", -- $0026d
          622 => x"84", -- $0026e
          623 => x"84", -- $0026f
          624 => x"84", -- $00270
          625 => x"85", -- $00271
          626 => x"85", -- $00272
          627 => x"85", -- $00273
          628 => x"85", -- $00274
          629 => x"85", -- $00275
          630 => x"85", -- $00276
          631 => x"85", -- $00277
          632 => x"85", -- $00278
          633 => x"85", -- $00279
          634 => x"85", -- $0027a
          635 => x"85", -- $0027b
          636 => x"85", -- $0027c
          637 => x"85", -- $0027d
          638 => x"85", -- $0027e
          639 => x"85", -- $0027f
          640 => x"85", -- $00280
          641 => x"85", -- $00281
          642 => x"85", -- $00282
          643 => x"85", -- $00283
          644 => x"85", -- $00284
          645 => x"85", -- $00285
          646 => x"85", -- $00286
          647 => x"85", -- $00287
          648 => x"85", -- $00288
          649 => x"85", -- $00289
          650 => x"85", -- $0028a
          651 => x"85", -- $0028b
          652 => x"85", -- $0028c
          653 => x"85", -- $0028d
          654 => x"85", -- $0028e
          655 => x"85", -- $0028f
          656 => x"85", -- $00290
          657 => x"85", -- $00291
          658 => x"85", -- $00292
          659 => x"86", -- $00293
          660 => x"85", -- $00294
          661 => x"85", -- $00295
          662 => x"86", -- $00296
          663 => x"86", -- $00297
          664 => x"86", -- $00298
          665 => x"86", -- $00299
          666 => x"86", -- $0029a
          667 => x"86", -- $0029b
          668 => x"86", -- $0029c
          669 => x"85", -- $0029d
          670 => x"85", -- $0029e
          671 => x"86", -- $0029f
          672 => x"86", -- $002a0
          673 => x"86", -- $002a1
          674 => x"86", -- $002a2
          675 => x"85", -- $002a3
          676 => x"86", -- $002a4
          677 => x"86", -- $002a5
          678 => x"86", -- $002a6
          679 => x"86", -- $002a7
          680 => x"86", -- $002a8
          681 => x"86", -- $002a9
          682 => x"85", -- $002aa
          683 => x"86", -- $002ab
          684 => x"85", -- $002ac
          685 => x"85", -- $002ad
          686 => x"86", -- $002ae
          687 => x"86", -- $002af
          688 => x"86", -- $002b0
          689 => x"86", -- $002b1
          690 => x"86", -- $002b2
          691 => x"86", -- $002b3
          692 => x"86", -- $002b4
          693 => x"86", -- $002b5
          694 => x"85", -- $002b6
          695 => x"85", -- $002b7
          696 => x"85", -- $002b8
          697 => x"85", -- $002b9
          698 => x"85", -- $002ba
          699 => x"85", -- $002bb
          700 => x"85", -- $002bc
          701 => x"85", -- $002bd
          702 => x"85", -- $002be
          703 => x"85", -- $002bf
          704 => x"85", -- $002c0
          705 => x"85", -- $002c1
          706 => x"85", -- $002c2
          707 => x"85", -- $002c3
          708 => x"85", -- $002c4
          709 => x"85", -- $002c5
          710 => x"84", -- $002c6
          711 => x"84", -- $002c7
          712 => x"85", -- $002c8
          713 => x"85", -- $002c9
          714 => x"85", -- $002ca
          715 => x"85", -- $002cb
          716 => x"85", -- $002cc
          717 => x"84", -- $002cd
          718 => x"84", -- $002ce
          719 => x"84", -- $002cf
          720 => x"84", -- $002d0
          721 => x"84", -- $002d1
          722 => x"84", -- $002d2
          723 => x"84", -- $002d3
          724 => x"84", -- $002d4
          725 => x"84", -- $002d5
          726 => x"84", -- $002d6
          727 => x"84", -- $002d7
          728 => x"84", -- $002d8
          729 => x"84", -- $002d9
          730 => x"84", -- $002da
          731 => x"84", -- $002db
          732 => x"84", -- $002dc
          733 => x"84", -- $002dd
          734 => x"83", -- $002de
          735 => x"83", -- $002df
          736 => x"83", -- $002e0
          737 => x"83", -- $002e1
          738 => x"83", -- $002e2
          739 => x"83", -- $002e3
          740 => x"83", -- $002e4
          741 => x"83", -- $002e5
          742 => x"83", -- $002e6
          743 => x"83", -- $002e7
          744 => x"83", -- $002e8
          745 => x"83", -- $002e9
          746 => x"83", -- $002ea
          747 => x"83", -- $002eb
          748 => x"83", -- $002ec
          749 => x"83", -- $002ed
          750 => x"83", -- $002ee
          751 => x"83", -- $002ef
          752 => x"83", -- $002f0
          753 => x"83", -- $002f1
          754 => x"83", -- $002f2
          755 => x"83", -- $002f3
          756 => x"83", -- $002f4
          757 => x"83", -- $002f5
          758 => x"83", -- $002f6
          759 => x"83", -- $002f7
          760 => x"82", -- $002f8
          761 => x"82", -- $002f9
          762 => x"82", -- $002fa
          763 => x"82", -- $002fb
          764 => x"82", -- $002fc
          765 => x"82", -- $002fd
          766 => x"82", -- $002fe
          767 => x"82", -- $002ff
          768 => x"82", -- $00300
          769 => x"83", -- $00301
          770 => x"82", -- $00302
          771 => x"82", -- $00303
          772 => x"82", -- $00304
          773 => x"82", -- $00305
          774 => x"82", -- $00306
          775 => x"82", -- $00307
          776 => x"82", -- $00308
          777 => x"82", -- $00309
          778 => x"82", -- $0030a
          779 => x"82", -- $0030b
          780 => x"82", -- $0030c
          781 => x"82", -- $0030d
          782 => x"82", -- $0030e
          783 => x"82", -- $0030f
          784 => x"82", -- $00310
          785 => x"82", -- $00311
          786 => x"82", -- $00312
          787 => x"82", -- $00313
          788 => x"82", -- $00314
          789 => x"82", -- $00315
          790 => x"82", -- $00316
          791 => x"82", -- $00317
          792 => x"82", -- $00318
          793 => x"82", -- $00319
          794 => x"82", -- $0031a
          795 => x"82", -- $0031b
          796 => x"82", -- $0031c
          797 => x"82", -- $0031d
          798 => x"82", -- $0031e
          799 => x"81", -- $0031f
          800 => x"81", -- $00320
          801 => x"81", -- $00321
          802 => x"81", -- $00322
          803 => x"81", -- $00323
          804 => x"81", -- $00324
          805 => x"81", -- $00325
          806 => x"81", -- $00326
          807 => x"81", -- $00327
          808 => x"81", -- $00328
          809 => x"81", -- $00329
          810 => x"81", -- $0032a
          811 => x"81", -- $0032b
          812 => x"81", -- $0032c
          813 => x"81", -- $0032d
          814 => x"81", -- $0032e
          815 => x"81", -- $0032f
          816 => x"81", -- $00330
          817 => x"81", -- $00331
          818 => x"80", -- $00332
          819 => x"81", -- $00333
          820 => x"81", -- $00334
          821 => x"81", -- $00335
          822 => x"81", -- $00336
          823 => x"81", -- $00337
          824 => x"81", -- $00338
          825 => x"80", -- $00339
          826 => x"80", -- $0033a
          827 => x"80", -- $0033b
          828 => x"80", -- $0033c
          829 => x"80", -- $0033d
          830 => x"80", -- $0033e
          831 => x"80", -- $0033f
          832 => x"80", -- $00340
          833 => x"80", -- $00341
          834 => x"80", -- $00342
          835 => x"80", -- $00343
          836 => x"80", -- $00344
          837 => x"80", -- $00345
          838 => x"80", -- $00346
          839 => x"80", -- $00347
          840 => x"80", -- $00348
          841 => x"80", -- $00349
          842 => x"80", -- $0034a
          843 => x"80", -- $0034b
          844 => x"80", -- $0034c
          845 => x"80", -- $0034d
          846 => x"80", -- $0034e
          847 => x"80", -- $0034f
          848 => x"80", -- $00350
          849 => x"80", -- $00351
          850 => x"80", -- $00352
          851 => x"80", -- $00353
          852 => x"80", -- $00354
          853 => x"80", -- $00355
          854 => x"80", -- $00356
          855 => x"7f", -- $00357
          856 => x"7f", -- $00358
          857 => x"80", -- $00359
          858 => x"80", -- $0035a
          859 => x"80", -- $0035b
          860 => x"80", -- $0035c
          861 => x"7f", -- $0035d
          862 => x"7f", -- $0035e
          863 => x"7f", -- $0035f
          864 => x"7f", -- $00360
          865 => x"7f", -- $00361
          866 => x"7f", -- $00362
          867 => x"7f", -- $00363
          868 => x"7f", -- $00364
          869 => x"7f", -- $00365
          870 => x"7f", -- $00366
          871 => x"7f", -- $00367
          872 => x"7f", -- $00368
          873 => x"7f", -- $00369
          874 => x"7f", -- $0036a
          875 => x"7e", -- $0036b
          876 => x"7e", -- $0036c
          877 => x"7e", -- $0036d
          878 => x"7e", -- $0036e
          879 => x"7e", -- $0036f
          880 => x"7e", -- $00370
          881 => x"7e", -- $00371
          882 => x"7e", -- $00372
          883 => x"7e", -- $00373
          884 => x"7e", -- $00374
          885 => x"7e", -- $00375
          886 => x"7e", -- $00376
          887 => x"7e", -- $00377
          888 => x"7e", -- $00378
          889 => x"7e", -- $00379
          890 => x"7e", -- $0037a
          891 => x"7e", -- $0037b
          892 => x"7e", -- $0037c
          893 => x"7e", -- $0037d
          894 => x"7e", -- $0037e
          895 => x"7e", -- $0037f
          896 => x"7e", -- $00380
          897 => x"7e", -- $00381
          898 => x"7e", -- $00382
          899 => x"7e", -- $00383
          900 => x"7e", -- $00384
          901 => x"7e", -- $00385
          902 => x"7e", -- $00386
          903 => x"7d", -- $00387
          904 => x"7d", -- $00388
          905 => x"7d", -- $00389
          906 => x"7d", -- $0038a
          907 => x"7d", -- $0038b
          908 => x"7d", -- $0038c
          909 => x"7d", -- $0038d
          910 => x"7d", -- $0038e
          911 => x"7d", -- $0038f
          912 => x"7d", -- $00390
          913 => x"7d", -- $00391
          914 => x"7d", -- $00392
          915 => x"7d", -- $00393
          916 => x"7d", -- $00394
          917 => x"7d", -- $00395
          918 => x"7d", -- $00396
          919 => x"7d", -- $00397
          920 => x"7d", -- $00398
          921 => x"7d", -- $00399
          922 => x"7d", -- $0039a
          923 => x"7d", -- $0039b
          924 => x"7d", -- $0039c
          925 => x"7d", -- $0039d
          926 => x"7d", -- $0039e
          927 => x"7d", -- $0039f
          928 => x"7d", -- $003a0
          929 => x"7d", -- $003a1
          930 => x"7d", -- $003a2
          931 => x"7d", -- $003a3
          932 => x"7d", -- $003a4
          933 => x"7d", -- $003a5
          934 => x"7d", -- $003a6
          935 => x"7d", -- $003a7
          936 => x"7d", -- $003a8
          937 => x"7d", -- $003a9
          938 => x"7d", -- $003aa
          939 => x"7d", -- $003ab
          940 => x"7d", -- $003ac
          941 => x"7d", -- $003ad
          942 => x"7d", -- $003ae
          943 => x"7d", -- $003af
          944 => x"7d", -- $003b0
          945 => x"7d", -- $003b1
          946 => x"7c", -- $003b2
          947 => x"7c", -- $003b3
          948 => x"7d", -- $003b4
          949 => x"7c", -- $003b5
          950 => x"7c", -- $003b6
          951 => x"7d", -- $003b7
          952 => x"7d", -- $003b8
          953 => x"7d", -- $003b9
          954 => x"7c", -- $003ba
          955 => x"7c", -- $003bb
          956 => x"7c", -- $003bc
          957 => x"7c", -- $003bd
          958 => x"7c", -- $003be
          959 => x"7c", -- $003bf
          960 => x"7c", -- $003c0
          961 => x"7c", -- $003c1
          962 => x"7c", -- $003c2
          963 => x"7c", -- $003c3
          964 => x"7c", -- $003c4
          965 => x"7c", -- $003c5
          966 => x"7c", -- $003c6
          967 => x"7c", -- $003c7
          968 => x"7c", -- $003c8
          969 => x"7c", -- $003c9
          970 => x"7c", -- $003ca
          971 => x"7c", -- $003cb
          972 => x"7c", -- $003cc
          973 => x"7c", -- $003cd
          974 => x"7c", -- $003ce
          975 => x"7c", -- $003cf
          976 => x"7c", -- $003d0
          977 => x"7c", -- $003d1
          978 => x"7c", -- $003d2
          979 => x"7c", -- $003d3
          980 => x"7c", -- $003d4
          981 => x"7c", -- $003d5
          982 => x"7c", -- $003d6
          983 => x"7c", -- $003d7
          984 => x"7c", -- $003d8
          985 => x"7b", -- $003d9
          986 => x"7b", -- $003da
          987 => x"7b", -- $003db
          988 => x"7b", -- $003dc
          989 => x"7b", -- $003dd
          990 => x"7c", -- $003de
          991 => x"7c", -- $003df
          992 => x"7c", -- $003e0
          993 => x"7c", -- $003e1
          994 => x"7b", -- $003e2
          995 => x"7b", -- $003e3
          996 => x"7b", -- $003e4
          997 => x"7b", -- $003e5
          998 => x"7b", -- $003e6
          999 => x"7b", -- $003e7
          1000 => x"7b", -- $003e8
          1001 => x"7b", -- $003e9
          1002 => x"7b", -- $003ea
          1003 => x"7b", -- $003eb
          1004 => x"7b", -- $003ec
          1005 => x"7b", -- $003ed
          1006 => x"7b", -- $003ee
          1007 => x"7b", -- $003ef
          1008 => x"7b", -- $003f0
          1009 => x"7b", -- $003f1
          1010 => x"7b", -- $003f2
          1011 => x"7b", -- $003f3
          1012 => x"7b", -- $003f4
          1013 => x"7b", -- $003f5
          1014 => x"7b", -- $003f6
          1015 => x"7b", -- $003f7
          1016 => x"7b", -- $003f8
          1017 => x"7b", -- $003f9
          1018 => x"7b", -- $003fa
          1019 => x"7b", -- $003fb
          1020 => x"7b", -- $003fc
          1021 => x"7a", -- $003fd
          1022 => x"7b", -- $003fe
          1023 => x"7b", -- $003ff
          1024 => x"7b", -- $00400
          1025 => x"7b", -- $00401
          1026 => x"7b", -- $00402
          1027 => x"7b", -- $00403
          1028 => x"7b", -- $00404
          1029 => x"7b", -- $00405
          1030 => x"7a", -- $00406
          1031 => x"7a", -- $00407
          1032 => x"7a", -- $00408
          1033 => x"7a", -- $00409
          1034 => x"7b", -- $0040a
          1035 => x"7b", -- $0040b
          1036 => x"7a", -- $0040c
          1037 => x"7a", -- $0040d
          1038 => x"7a", -- $0040e
          1039 => x"7a", -- $0040f
          1040 => x"7a", -- $00410
          1041 => x"7b", -- $00411
          1042 => x"7b", -- $00412
          1043 => x"7b", -- $00413
          1044 => x"7b", -- $00414
          1045 => x"7b", -- $00415
          1046 => x"7a", -- $00416
          1047 => x"7a", -- $00417
          1048 => x"7a", -- $00418
          1049 => x"7a", -- $00419
          1050 => x"7a", -- $0041a
          1051 => x"7a", -- $0041b
          1052 => x"7a", -- $0041c
          1053 => x"7b", -- $0041d
          1054 => x"7b", -- $0041e
          1055 => x"7b", -- $0041f
          1056 => x"7b", -- $00420
          1057 => x"7b", -- $00421
          1058 => x"7b", -- $00422
          1059 => x"7b", -- $00423
          1060 => x"7b", -- $00424
          1061 => x"7b", -- $00425
          1062 => x"7b", -- $00426
          1063 => x"7b", -- $00427
          1064 => x"7b", -- $00428
          1065 => x"7b", -- $00429
          1066 => x"7b", -- $0042a
          1067 => x"7b", -- $0042b
          1068 => x"7b", -- $0042c
          1069 => x"7b", -- $0042d
          1070 => x"7b", -- $0042e
          1071 => x"7b", -- $0042f
          1072 => x"7b", -- $00430
          1073 => x"7b", -- $00431
          1074 => x"7b", -- $00432
          1075 => x"7b", -- $00433
          1076 => x"7b", -- $00434
          1077 => x"7b", -- $00435
          1078 => x"7b", -- $00436
          1079 => x"7b", -- $00437
          1080 => x"7b", -- $00438
          1081 => x"7b", -- $00439
          1082 => x"7b", -- $0043a
          1083 => x"7b", -- $0043b
          1084 => x"7c", -- $0043c
          1085 => x"7c", -- $0043d
          1086 => x"7c", -- $0043e
          1087 => x"7c", -- $0043f
          1088 => x"7c", -- $00440
          1089 => x"7c", -- $00441
          1090 => x"7c", -- $00442
          1091 => x"7c", -- $00443
          1092 => x"7c", -- $00444
          1093 => x"7c", -- $00445
          1094 => x"7c", -- $00446
          1095 => x"7c", -- $00447
          1096 => x"7c", -- $00448
          1097 => x"7c", -- $00449
          1098 => x"7c", -- $0044a
          1099 => x"7c", -- $0044b
          1100 => x"7c", -- $0044c
          1101 => x"7c", -- $0044d
          1102 => x"7c", -- $0044e
          1103 => x"7c", -- $0044f
          1104 => x"7c", -- $00450
          1105 => x"7c", -- $00451
          1106 => x"7d", -- $00452
          1107 => x"7d", -- $00453
          1108 => x"7d", -- $00454
          1109 => x"7d", -- $00455
          1110 => x"7d", -- $00456
          1111 => x"7d", -- $00457
          1112 => x"7d", -- $00458
          1113 => x"7d", -- $00459
          1114 => x"7d", -- $0045a
          1115 => x"7d", -- $0045b
          1116 => x"7d", -- $0045c
          1117 => x"7d", -- $0045d
          1118 => x"7d", -- $0045e
          1119 => x"7d", -- $0045f
          1120 => x"7d", -- $00460
          1121 => x"7d", -- $00461
          1122 => x"7d", -- $00462
          1123 => x"7d", -- $00463
          1124 => x"7d", -- $00464
          1125 => x"7d", -- $00465
          1126 => x"7d", -- $00466
          1127 => x"7d", -- $00467
          1128 => x"7d", -- $00468
          1129 => x"7d", -- $00469
          1130 => x"7d", -- $0046a
          1131 => x"7d", -- $0046b
          1132 => x"7d", -- $0046c
          1133 => x"7d", -- $0046d
          1134 => x"7d", -- $0046e
          1135 => x"7d", -- $0046f
          1136 => x"7d", -- $00470
          1137 => x"7e", -- $00471
          1138 => x"7d", -- $00472
          1139 => x"7d", -- $00473
          1140 => x"7d", -- $00474
          1141 => x"7d", -- $00475
          1142 => x"7d", -- $00476
          1143 => x"7d", -- $00477
          1144 => x"7e", -- $00478
          1145 => x"7e", -- $00479
          1146 => x"7e", -- $0047a
          1147 => x"7e", -- $0047b
          1148 => x"7d", -- $0047c
          1149 => x"7e", -- $0047d
          1150 => x"7e", -- $0047e
          1151 => x"7e", -- $0047f
          1152 => x"7e", -- $00480
          1153 => x"7e", -- $00481
          1154 => x"7e", -- $00482
          1155 => x"7e", -- $00483
          1156 => x"7e", -- $00484
          1157 => x"7e", -- $00485
          1158 => x"7e", -- $00486
          1159 => x"7e", -- $00487
          1160 => x"7e", -- $00488
          1161 => x"7e", -- $00489
          1162 => x"7e", -- $0048a
          1163 => x"7e", -- $0048b
          1164 => x"7e", -- $0048c
          1165 => x"7e", -- $0048d
          1166 => x"7e", -- $0048e
          1167 => x"7e", -- $0048f
          1168 => x"7e", -- $00490
          1169 => x"7e", -- $00491
          1170 => x"7e", -- $00492
          1171 => x"7e", -- $00493
          1172 => x"7e", -- $00494
          1173 => x"7e", -- $00495
          1174 => x"7e", -- $00496
          1175 => x"7e", -- $00497
          1176 => x"7e", -- $00498
          1177 => x"7e", -- $00499
          1178 => x"7e", -- $0049a
          1179 => x"7e", -- $0049b
          1180 => x"7e", -- $0049c
          1181 => x"7e", -- $0049d
          1182 => x"7e", -- $0049e
          1183 => x"7e", -- $0049f
          1184 => x"7e", -- $004a0
          1185 => x"7e", -- $004a1
          1186 => x"7e", -- $004a2
          1187 => x"7e", -- $004a3
          1188 => x"7e", -- $004a4
          1189 => x"7e", -- $004a5
          1190 => x"7e", -- $004a6
          1191 => x"7e", -- $004a7
          1192 => x"7e", -- $004a8
          1193 => x"7e", -- $004a9
          1194 => x"7e", -- $004aa
          1195 => x"7f", -- $004ab
          1196 => x"7f", -- $004ac
          1197 => x"7f", -- $004ad
          1198 => x"7f", -- $004ae
          1199 => x"7f", -- $004af
          1200 => x"7f", -- $004b0
          1201 => x"7f", -- $004b1
          1202 => x"7f", -- $004b2
          1203 => x"7f", -- $004b3
          1204 => x"7f", -- $004b4
          1205 => x"7f", -- $004b5
          1206 => x"7f", -- $004b6
          1207 => x"7f", -- $004b7
          1208 => x"7f", -- $004b8
          1209 => x"7f", -- $004b9
          1210 => x"7f", -- $004ba
          1211 => x"7f", -- $004bb
          1212 => x"7f", -- $004bc
          1213 => x"7f", -- $004bd
          1214 => x"7f", -- $004be
          1215 => x"7f", -- $004bf
          1216 => x"7f", -- $004c0
          1217 => x"7f", -- $004c1
          1218 => x"80", -- $004c2
          1219 => x"80", -- $004c3
          1220 => x"80", -- $004c4
          1221 => x"80", -- $004c5
          1222 => x"80", -- $004c6
          1223 => x"80", -- $004c7
          1224 => x"80", -- $004c8
          1225 => x"80", -- $004c9
          1226 => x"80", -- $004ca
          1227 => x"80", -- $004cb
          1228 => x"80", -- $004cc
          1229 => x"80", -- $004cd
          1230 => x"80", -- $004ce
          1231 => x"80", -- $004cf
          1232 => x"80", -- $004d0
          1233 => x"80", -- $004d1
          1234 => x"80", -- $004d2
          1235 => x"80", -- $004d3
          1236 => x"80", -- $004d4
          1237 => x"80", -- $004d5
          1238 => x"80", -- $004d6
          1239 => x"80", -- $004d7
          1240 => x"80", -- $004d8
          1241 => x"80", -- $004d9
          1242 => x"80", -- $004da
          1243 => x"80", -- $004db
          1244 => x"80", -- $004dc
          1245 => x"80", -- $004dd
          1246 => x"80", -- $004de
          1247 => x"80", -- $004df
          1248 => x"80", -- $004e0
          1249 => x"80", -- $004e1
          1250 => x"80", -- $004e2
          1251 => x"80", -- $004e3
          1252 => x"80", -- $004e4
          1253 => x"80", -- $004e5
          1254 => x"80", -- $004e6
          1255 => x"80", -- $004e7
          1256 => x"80", -- $004e8
          1257 => x"80", -- $004e9
          1258 => x"81", -- $004ea
          1259 => x"80", -- $004eb
          1260 => x"81", -- $004ec
          1261 => x"81", -- $004ed
          1262 => x"81", -- $004ee
          1263 => x"81", -- $004ef
          1264 => x"81", -- $004f0
          1265 => x"81", -- $004f1
          1266 => x"81", -- $004f2
          1267 => x"81", -- $004f3
          1268 => x"81", -- $004f4
          1269 => x"81", -- $004f5
          1270 => x"81", -- $004f6
          1271 => x"81", -- $004f7
          1272 => x"81", -- $004f8
          1273 => x"81", -- $004f9
          1274 => x"81", -- $004fa
          1275 => x"81", -- $004fb
          1276 => x"81", -- $004fc
          1277 => x"81", -- $004fd
          1278 => x"81", -- $004fe
          1279 => x"81", -- $004ff
          1280 => x"81", -- $00500
          1281 => x"81", -- $00501
          1282 => x"81", -- $00502
          1283 => x"81", -- $00503
          1284 => x"81", -- $00504
          1285 => x"81", -- $00505
          1286 => x"81", -- $00506
          1287 => x"81", -- $00507
          1288 => x"82", -- $00508
          1289 => x"82", -- $00509
          1290 => x"82", -- $0050a
          1291 => x"82", -- $0050b
          1292 => x"82", -- $0050c
          1293 => x"82", -- $0050d
          1294 => x"82", -- $0050e
          1295 => x"82", -- $0050f
          1296 => x"82", -- $00510
          1297 => x"82", -- $00511
          1298 => x"82", -- $00512
          1299 => x"82", -- $00513
          1300 => x"82", -- $00514
          1301 => x"82", -- $00515
          1302 => x"82", -- $00516
          1303 => x"83", -- $00517
          1304 => x"83", -- $00518
          1305 => x"83", -- $00519
          1306 => x"82", -- $0051a
          1307 => x"82", -- $0051b
          1308 => x"83", -- $0051c
          1309 => x"83", -- $0051d
          1310 => x"82", -- $0051e
          1311 => x"82", -- $0051f
          1312 => x"82", -- $00520
          1313 => x"83", -- $00521
          1314 => x"83", -- $00522
          1315 => x"83", -- $00523
          1316 => x"83", -- $00524
          1317 => x"83", -- $00525
          1318 => x"83", -- $00526
          1319 => x"83", -- $00527
          1320 => x"83", -- $00528
          1321 => x"83", -- $00529
          1322 => x"83", -- $0052a
          1323 => x"83", -- $0052b
          1324 => x"83", -- $0052c
          1325 => x"83", -- $0052d
          1326 => x"83", -- $0052e
          1327 => x"83", -- $0052f
          1328 => x"83", -- $00530
          1329 => x"83", -- $00531
          1330 => x"83", -- $00532
          1331 => x"83", -- $00533
          1332 => x"83", -- $00534
          1333 => x"83", -- $00535
          1334 => x"83", -- $00536
          1335 => x"84", -- $00537
          1336 => x"83", -- $00538
          1337 => x"83", -- $00539
          1338 => x"83", -- $0053a
          1339 => x"83", -- $0053b
          1340 => x"83", -- $0053c
          1341 => x"83", -- $0053d
          1342 => x"84", -- $0053e
          1343 => x"84", -- $0053f
          1344 => x"84", -- $00540
          1345 => x"84", -- $00541
          1346 => x"83", -- $00542
          1347 => x"83", -- $00543
          1348 => x"83", -- $00544
          1349 => x"83", -- $00545
          1350 => x"83", -- $00546
          1351 => x"83", -- $00547
          1352 => x"84", -- $00548
          1353 => x"84", -- $00549
          1354 => x"84", -- $0054a
          1355 => x"84", -- $0054b
          1356 => x"83", -- $0054c
          1357 => x"83", -- $0054d
          1358 => x"83", -- $0054e
          1359 => x"84", -- $0054f
          1360 => x"84", -- $00550
          1361 => x"84", -- $00551
          1362 => x"84", -- $00552
          1363 => x"83", -- $00553
          1364 => x"83", -- $00554
          1365 => x"84", -- $00555
          1366 => x"84", -- $00556
          1367 => x"84", -- $00557
          1368 => x"84", -- $00558
          1369 => x"84", -- $00559
          1370 => x"84", -- $0055a
          1371 => x"84", -- $0055b
          1372 => x"84", -- $0055c
          1373 => x"84", -- $0055d
          1374 => x"84", -- $0055e
          1375 => x"84", -- $0055f
          1376 => x"84", -- $00560
          1377 => x"84", -- $00561
          1378 => x"84", -- $00562
          1379 => x"84", -- $00563
          1380 => x"84", -- $00564
          1381 => x"84", -- $00565
          1382 => x"84", -- $00566
          1383 => x"84", -- $00567
          1384 => x"84", -- $00568
          1385 => x"84", -- $00569
          1386 => x"84", -- $0056a
          1387 => x"84", -- $0056b
          1388 => x"84", -- $0056c
          1389 => x"84", -- $0056d
          1390 => x"84", -- $0056e
          1391 => x"84", -- $0056f
          1392 => x"84", -- $00570
          1393 => x"85", -- $00571
          1394 => x"85", -- $00572
          1395 => x"85", -- $00573
          1396 => x"85", -- $00574
          1397 => x"85", -- $00575
          1398 => x"85", -- $00576
          1399 => x"85", -- $00577
          1400 => x"85", -- $00578
          1401 => x"85", -- $00579
          1402 => x"85", -- $0057a
          1403 => x"85", -- $0057b
          1404 => x"85", -- $0057c
          1405 => x"85", -- $0057d
          1406 => x"85", -- $0057e
          1407 => x"85", -- $0057f
          1408 => x"85", -- $00580
          1409 => x"85", -- $00581
          1410 => x"85", -- $00582
          1411 => x"85", -- $00583
          1412 => x"85", -- $00584
          1413 => x"85", -- $00585
          1414 => x"85", -- $00586
          1415 => x"85", -- $00587
          1416 => x"85", -- $00588
          1417 => x"85", -- $00589
          1418 => x"85", -- $0058a
          1419 => x"85", -- $0058b
          1420 => x"85", -- $0058c
          1421 => x"85", -- $0058d
          1422 => x"85", -- $0058e
          1423 => x"85", -- $0058f
          1424 => x"85", -- $00590
          1425 => x"85", -- $00591
          1426 => x"85", -- $00592
          1427 => x"85", -- $00593
          1428 => x"85", -- $00594
          1429 => x"85", -- $00595
          1430 => x"85", -- $00596
          1431 => x"85", -- $00597
          1432 => x"85", -- $00598
          1433 => x"85", -- $00599
          1434 => x"84", -- $0059a
          1435 => x"84", -- $0059b
          1436 => x"85", -- $0059c
          1437 => x"85", -- $0059d
          1438 => x"85", -- $0059e
          1439 => x"84", -- $0059f
          1440 => x"84", -- $005a0
          1441 => x"84", -- $005a1
          1442 => x"84", -- $005a2
          1443 => x"84", -- $005a3
          1444 => x"84", -- $005a4
          1445 => x"84", -- $005a5
          1446 => x"84", -- $005a6
          1447 => x"84", -- $005a7
          1448 => x"84", -- $005a8
          1449 => x"84", -- $005a9
          1450 => x"84", -- $005aa
          1451 => x"84", -- $005ab
          1452 => x"84", -- $005ac
          1453 => x"84", -- $005ad
          1454 => x"84", -- $005ae
          1455 => x"84", -- $005af
          1456 => x"84", -- $005b0
          1457 => x"84", -- $005b1
          1458 => x"85", -- $005b2
          1459 => x"84", -- $005b3
          1460 => x"85", -- $005b4
          1461 => x"85", -- $005b5
          1462 => x"85", -- $005b6
          1463 => x"85", -- $005b7
          1464 => x"85", -- $005b8
          1465 => x"84", -- $005b9
          1466 => x"84", -- $005ba
          1467 => x"84", -- $005bb
          1468 => x"84", -- $005bc
          1469 => x"84", -- $005bd
          1470 => x"84", -- $005be
          1471 => x"84", -- $005bf
          1472 => x"84", -- $005c0
          1473 => x"84", -- $005c1
          1474 => x"84", -- $005c2
          1475 => x"84", -- $005c3
          1476 => x"84", -- $005c4
          1477 => x"84", -- $005c5
          1478 => x"84", -- $005c6
          1479 => x"84", -- $005c7
          1480 => x"84", -- $005c8
          1481 => x"84", -- $005c9
          1482 => x"84", -- $005ca
          1483 => x"84", -- $005cb
          1484 => x"84", -- $005cc
          1485 => x"84", -- $005cd
          1486 => x"84", -- $005ce
          1487 => x"84", -- $005cf
          1488 => x"84", -- $005d0
          1489 => x"84", -- $005d1
          1490 => x"84", -- $005d2
          1491 => x"84", -- $005d3
          1492 => x"84", -- $005d4
          1493 => x"84", -- $005d5
          1494 => x"84", -- $005d6
          1495 => x"84", -- $005d7
          1496 => x"84", -- $005d8
          1497 => x"84", -- $005d9
          1498 => x"84", -- $005da
          1499 => x"84", -- $005db
          1500 => x"84", -- $005dc
          1501 => x"84", -- $005dd
          1502 => x"84", -- $005de
          1503 => x"84", -- $005df
          1504 => x"84", -- $005e0
          1505 => x"84", -- $005e1
          1506 => x"84", -- $005e2
          1507 => x"84", -- $005e3
          1508 => x"84", -- $005e4
          1509 => x"84", -- $005e5
          1510 => x"84", -- $005e6
          1511 => x"84", -- $005e7
          1512 => x"84", -- $005e8
          1513 => x"84", -- $005e9
          1514 => x"84", -- $005ea
          1515 => x"84", -- $005eb
          1516 => x"84", -- $005ec
          1517 => x"84", -- $005ed
          1518 => x"83", -- $005ee
          1519 => x"83", -- $005ef
          1520 => x"83", -- $005f0
          1521 => x"83", -- $005f1
          1522 => x"83", -- $005f2
          1523 => x"83", -- $005f3
          1524 => x"84", -- $005f4
          1525 => x"83", -- $005f5
          1526 => x"83", -- $005f6
          1527 => x"83", -- $005f7
          1528 => x"83", -- $005f8
          1529 => x"83", -- $005f9
          1530 => x"83", -- $005fa
          1531 => x"83", -- $005fb
          1532 => x"83", -- $005fc
          1533 => x"83", -- $005fd
          1534 => x"83", -- $005fe
          1535 => x"83", -- $005ff
          1536 => x"83", -- $00600
          1537 => x"83", -- $00601
          1538 => x"83", -- $00602
          1539 => x"83", -- $00603
          1540 => x"83", -- $00604
          1541 => x"83", -- $00605
          1542 => x"82", -- $00606
          1543 => x"82", -- $00607
          1544 => x"82", -- $00608
          1545 => x"82", -- $00609
          1546 => x"82", -- $0060a
          1547 => x"82", -- $0060b
          1548 => x"82", -- $0060c
          1549 => x"82", -- $0060d
          1550 => x"82", -- $0060e
          1551 => x"82", -- $0060f
          1552 => x"82", -- $00610
          1553 => x"82", -- $00611
          1554 => x"82", -- $00612
          1555 => x"82", -- $00613
          1556 => x"82", -- $00614
          1557 => x"82", -- $00615
          1558 => x"82", -- $00616
          1559 => x"82", -- $00617
          1560 => x"82", -- $00618
          1561 => x"82", -- $00619
          1562 => x"82", -- $0061a
          1563 => x"81", -- $0061b
          1564 => x"81", -- $0061c
          1565 => x"81", -- $0061d
          1566 => x"81", -- $0061e
          1567 => x"81", -- $0061f
          1568 => x"81", -- $00620
          1569 => x"81", -- $00621
          1570 => x"81", -- $00622
          1571 => x"81", -- $00623
          1572 => x"81", -- $00624
          1573 => x"81", -- $00625
          1574 => x"81", -- $00626
          1575 => x"81", -- $00627
          1576 => x"81", -- $00628
          1577 => x"81", -- $00629
          1578 => x"81", -- $0062a
          1579 => x"81", -- $0062b
          1580 => x"81", -- $0062c
          1581 => x"81", -- $0062d
          1582 => x"81", -- $0062e
          1583 => x"81", -- $0062f
          1584 => x"81", -- $00630
          1585 => x"81", -- $00631
          1586 => x"81", -- $00632
          1587 => x"81", -- $00633
          1588 => x"81", -- $00634
          1589 => x"81", -- $00635
          1590 => x"81", -- $00636
          1591 => x"80", -- $00637
          1592 => x"81", -- $00638
          1593 => x"81", -- $00639
          1594 => x"81", -- $0063a
          1595 => x"80", -- $0063b
          1596 => x"80", -- $0063c
          1597 => x"80", -- $0063d
          1598 => x"80", -- $0063e
          1599 => x"80", -- $0063f
          1600 => x"80", -- $00640
          1601 => x"81", -- $00641
          1602 => x"80", -- $00642
          1603 => x"80", -- $00643
          1604 => x"80", -- $00644
          1605 => x"80", -- $00645
          1606 => x"80", -- $00646
          1607 => x"80", -- $00647
          1608 => x"80", -- $00648
          1609 => x"80", -- $00649
          1610 => x"80", -- $0064a
          1611 => x"80", -- $0064b
          1612 => x"80", -- $0064c
          1613 => x"80", -- $0064d
          1614 => x"80", -- $0064e
          1615 => x"80", -- $0064f
          1616 => x"80", -- $00650
          1617 => x"80", -- $00651
          1618 => x"80", -- $00652
          1619 => x"80", -- $00653
          1620 => x"80", -- $00654
          1621 => x"80", -- $00655
          1622 => x"80", -- $00656
          1623 => x"80", -- $00657
          1624 => x"80", -- $00658
          1625 => x"80", -- $00659
          1626 => x"80", -- $0065a
          1627 => x"80", -- $0065b
          1628 => x"80", -- $0065c
          1629 => x"80", -- $0065d
          1630 => x"80", -- $0065e
          1631 => x"80", -- $0065f
          1632 => x"80", -- $00660
          1633 => x"80", -- $00661
          1634 => x"7f", -- $00662
          1635 => x"7f", -- $00663
          1636 => x"7f", -- $00664
          1637 => x"7f", -- $00665
          1638 => x"7f", -- $00666
          1639 => x"7f", -- $00667
          1640 => x"7f", -- $00668
          1641 => x"7f", -- $00669
          1642 => x"7f", -- $0066a
          1643 => x"7f", -- $0066b
          1644 => x"7f", -- $0066c
          1645 => x"7f", -- $0066d
          1646 => x"7f", -- $0066e
          1647 => x"7f", -- $0066f
          1648 => x"7f", -- $00670
          1649 => x"7f", -- $00671
          1650 => x"7f", -- $00672
          1651 => x"7e", -- $00673
          1652 => x"7f", -- $00674
          1653 => x"7f", -- $00675
          1654 => x"7f", -- $00676
          1655 => x"7e", -- $00677
          1656 => x"7e", -- $00678
          1657 => x"7e", -- $00679
          1658 => x"7e", -- $0067a
          1659 => x"7e", -- $0067b
          1660 => x"7e", -- $0067c
          1661 => x"7e", -- $0067d
          1662 => x"7e", -- $0067e
          1663 => x"7e", -- $0067f
          1664 => x"7e", -- $00680
          1665 => x"7e", -- $00681
          1666 => x"7e", -- $00682
          1667 => x"7e", -- $00683
          1668 => x"7e", -- $00684
          1669 => x"7e", -- $00685
          1670 => x"7e", -- $00686
          1671 => x"7e", -- $00687
          1672 => x"7d", -- $00688
          1673 => x"7d", -- $00689
          1674 => x"7d", -- $0068a
          1675 => x"7d", -- $0068b
          1676 => x"7d", -- $0068c
          1677 => x"7d", -- $0068d
          1678 => x"7d", -- $0068e
          1679 => x"7d", -- $0068f
          1680 => x"7d", -- $00690
          1681 => x"7d", -- $00691
          1682 => x"7d", -- $00692
          1683 => x"7d", -- $00693
          1684 => x"7d", -- $00694
          1685 => x"7d", -- $00695
          1686 => x"7d", -- $00696
          1687 => x"7d", -- $00697
          1688 => x"7d", -- $00698
          1689 => x"7d", -- $00699
          1690 => x"7d", -- $0069a
          1691 => x"7d", -- $0069b
          1692 => x"7d", -- $0069c
          1693 => x"7d", -- $0069d
          1694 => x"7d", -- $0069e
          1695 => x"7d", -- $0069f
          1696 => x"7d", -- $006a0
          1697 => x"7d", -- $006a1
          1698 => x"7d", -- $006a2
          1699 => x"7d", -- $006a3
          1700 => x"7d", -- $006a4
          1701 => x"7d", -- $006a5
          1702 => x"7d", -- $006a6
          1703 => x"7d", -- $006a7
          1704 => x"7d", -- $006a8
          1705 => x"7d", -- $006a9
          1706 => x"7d", -- $006aa
          1707 => x"7d", -- $006ab
          1708 => x"7d", -- $006ac
          1709 => x"7d", -- $006ad
          1710 => x"7d", -- $006ae
          1711 => x"7d", -- $006af
          1712 => x"7d", -- $006b0
          1713 => x"7d", -- $006b1
          1714 => x"7d", -- $006b2
          1715 => x"7c", -- $006b3
          1716 => x"7d", -- $006b4
          1717 => x"7d", -- $006b5
          1718 => x"7d", -- $006b6
          1719 => x"7d", -- $006b7
          1720 => x"7d", -- $006b8
          1721 => x"7d", -- $006b9
          1722 => x"7d", -- $006ba
          1723 => x"7d", -- $006bb
          1724 => x"7d", -- $006bc
          1725 => x"7d", -- $006bd
          1726 => x"7d", -- $006be
          1727 => x"7d", -- $006bf
          1728 => x"7d", -- $006c0
          1729 => x"7d", -- $006c1
          1730 => x"7d", -- $006c2
          1731 => x"7d", -- $006c3
          1732 => x"7d", -- $006c4
          1733 => x"7d", -- $006c5
          1734 => x"7d", -- $006c6
          1735 => x"7d", -- $006c7
          1736 => x"7d", -- $006c8
          1737 => x"7d", -- $006c9
          1738 => x"7d", -- $006ca
          1739 => x"7d", -- $006cb
          1740 => x"7d", -- $006cc
          1741 => x"7d", -- $006cd
          1742 => x"7d", -- $006ce
          1743 => x"7d", -- $006cf
          1744 => x"7d", -- $006d0
          1745 => x"7d", -- $006d1
          1746 => x"7d", -- $006d2
          1747 => x"7d", -- $006d3
          1748 => x"7d", -- $006d4
          1749 => x"7d", -- $006d5
          1750 => x"7d", -- $006d6
          1751 => x"7d", -- $006d7
          1752 => x"7d", -- $006d8
          1753 => x"7d", -- $006d9
          1754 => x"7d", -- $006da
          1755 => x"7d", -- $006db
          1756 => x"7d", -- $006dc
          1757 => x"7d", -- $006dd
          1758 => x"7d", -- $006de
          1759 => x"7d", -- $006df
          1760 => x"7d", -- $006e0
          1761 => x"7d", -- $006e1
          1762 => x"7d", -- $006e2
          1763 => x"7d", -- $006e3
          1764 => x"7d", -- $006e4
          1765 => x"7d", -- $006e5
          1766 => x"7d", -- $006e6
          1767 => x"7d", -- $006e7
          1768 => x"7d", -- $006e8
          1769 => x"7d", -- $006e9
          1770 => x"7d", -- $006ea
          1771 => x"7d", -- $006eb
          1772 => x"7d", -- $006ec
          1773 => x"7d", -- $006ed
          1774 => x"7d", -- $006ee
          1775 => x"7d", -- $006ef
          1776 => x"7d", -- $006f0
          1777 => x"7d", -- $006f1
          1778 => x"7d", -- $006f2
          1779 => x"7d", -- $006f3
          1780 => x"7d", -- $006f4
          1781 => x"7d", -- $006f5
          1782 => x"7d", -- $006f6
          1783 => x"7d", -- $006f7
          1784 => x"7d", -- $006f8
          1785 => x"7d", -- $006f9
          1786 => x"7c", -- $006fa
          1787 => x"7c", -- $006fb
          1788 => x"7c", -- $006fc
          1789 => x"7c", -- $006fd
          1790 => x"7c", -- $006fe
          1791 => x"7c", -- $006ff
          1792 => x"7c", -- $00700
          1793 => x"7c", -- $00701
          1794 => x"7c", -- $00702
          1795 => x"7c", -- $00703
          1796 => x"7c", -- $00704
          1797 => x"7c", -- $00705
          1798 => x"7c", -- $00706
          1799 => x"7c", -- $00707
          1800 => x"7c", -- $00708
          1801 => x"7c", -- $00709
          1802 => x"7c", -- $0070a
          1803 => x"7c", -- $0070b
          1804 => x"7c", -- $0070c
          1805 => x"7c", -- $0070d
          1806 => x"7c", -- $0070e
          1807 => x"7c", -- $0070f
          1808 => x"7c", -- $00710
          1809 => x"7c", -- $00711
          1810 => x"7c", -- $00712
          1811 => x"7c", -- $00713
          1812 => x"7c", -- $00714
          1813 => x"7c", -- $00715
          1814 => x"7c", -- $00716
          1815 => x"7c", -- $00717
          1816 => x"7c", -- $00718
          1817 => x"7c", -- $00719
          1818 => x"7c", -- $0071a
          1819 => x"7c", -- $0071b
          1820 => x"7c", -- $0071c
          1821 => x"7c", -- $0071d
          1822 => x"7c", -- $0071e
          1823 => x"7c", -- $0071f
          1824 => x"7c", -- $00720
          1825 => x"7c", -- $00721
          1826 => x"7c", -- $00722
          1827 => x"7b", -- $00723
          1828 => x"7b", -- $00724
          1829 => x"7b", -- $00725
          1830 => x"7b", -- $00726
          1831 => x"7b", -- $00727
          1832 => x"7b", -- $00728
          1833 => x"7b", -- $00729
          1834 => x"7b", -- $0072a
          1835 => x"7b", -- $0072b
          1836 => x"7c", -- $0072c
          1837 => x"7c", -- $0072d
          1838 => x"7c", -- $0072e
          1839 => x"7b", -- $0072f
          1840 => x"7b", -- $00730
          1841 => x"7b", -- $00731
          1842 => x"7b", -- $00732
          1843 => x"7b", -- $00733
          1844 => x"7c", -- $00734
          1845 => x"7b", -- $00735
          1846 => x"7b", -- $00736
          1847 => x"7b", -- $00737
          1848 => x"7b", -- $00738
          1849 => x"7b", -- $00739
          1850 => x"7b", -- $0073a
          1851 => x"7b", -- $0073b
          1852 => x"7b", -- $0073c
          1853 => x"7b", -- $0073d
          1854 => x"7b", -- $0073e
          1855 => x"7b", -- $0073f
          1856 => x"7b", -- $00740
          1857 => x"7b", -- $00741
          1858 => x"7b", -- $00742
          1859 => x"7b", -- $00743
          1860 => x"7b", -- $00744
          1861 => x"7b", -- $00745
          1862 => x"7b", -- $00746
          1863 => x"7b", -- $00747
          1864 => x"7b", -- $00748
          1865 => x"7b", -- $00749
          1866 => x"7b", -- $0074a
          1867 => x"7b", -- $0074b
          1868 => x"7c", -- $0074c
          1869 => x"7b", -- $0074d
          1870 => x"7b", -- $0074e
          1871 => x"7b", -- $0074f
          1872 => x"7b", -- $00750
          1873 => x"7b", -- $00751
          1874 => x"7b", -- $00752
          1875 => x"7b", -- $00753
          1876 => x"7b", -- $00754
          1877 => x"7c", -- $00755
          1878 => x"7c", -- $00756
          1879 => x"7c", -- $00757
          1880 => x"7c", -- $00758
          1881 => x"7b", -- $00759
          1882 => x"7b", -- $0075a
          1883 => x"7c", -- $0075b
          1884 => x"7c", -- $0075c
          1885 => x"7c", -- $0075d
          1886 => x"7c", -- $0075e
          1887 => x"7c", -- $0075f
          1888 => x"7c", -- $00760
          1889 => x"7c", -- $00761
          1890 => x"7c", -- $00762
          1891 => x"7c", -- $00763
          1892 => x"7c", -- $00764
          1893 => x"7c", -- $00765
          1894 => x"7c", -- $00766
          1895 => x"7c", -- $00767
          1896 => x"7d", -- $00768
          1897 => x"7d", -- $00769
          1898 => x"7d", -- $0076a
          1899 => x"7c", -- $0076b
          1900 => x"7c", -- $0076c
          1901 => x"7c", -- $0076d
          1902 => x"7d", -- $0076e
          1903 => x"7d", -- $0076f
          1904 => x"7d", -- $00770
          1905 => x"7d", -- $00771
          1906 => x"7d", -- $00772
          1907 => x"7d", -- $00773
          1908 => x"7d", -- $00774
          1909 => x"7d", -- $00775
          1910 => x"7e", -- $00776
          1911 => x"7d", -- $00777
          1912 => x"7d", -- $00778
          1913 => x"7d", -- $00779
          1914 => x"7d", -- $0077a
          1915 => x"7d", -- $0077b
          1916 => x"7e", -- $0077c
          1917 => x"7e", -- $0077d
          1918 => x"7d", -- $0077e
          1919 => x"7d", -- $0077f
          1920 => x"7e", -- $00780
          1921 => x"7e", -- $00781
          1922 => x"7e", -- $00782
          1923 => x"7e", -- $00783
          1924 => x"7e", -- $00784
          1925 => x"7e", -- $00785
          1926 => x"7e", -- $00786
          1927 => x"7e", -- $00787
          1928 => x"7f", -- $00788
          1929 => x"7f", -- $00789
          1930 => x"7f", -- $0078a
          1931 => x"7e", -- $0078b
          1932 => x"7e", -- $0078c
          1933 => x"7e", -- $0078d
          1934 => x"7e", -- $0078e
          1935 => x"7f", -- $0078f
          1936 => x"7f", -- $00790
          1937 => x"7f", -- $00791
          1938 => x"7f", -- $00792
          1939 => x"7f", -- $00793
          1940 => x"7f", -- $00794
          1941 => x"7f", -- $00795
          1942 => x"7f", -- $00796
          1943 => x"7f", -- $00797
          1944 => x"7f", -- $00798
          1945 => x"7f", -- $00799
          1946 => x"7f", -- $0079a
          1947 => x"7f", -- $0079b
          1948 => x"7f", -- $0079c
          1949 => x"7f", -- $0079d
          1950 => x"7f", -- $0079e
          1951 => x"7f", -- $0079f
          1952 => x"7f", -- $007a0
          1953 => x"80", -- $007a1
          1954 => x"80", -- $007a2
          1955 => x"80", -- $007a3
          1956 => x"7f", -- $007a4
          1957 => x"7f", -- $007a5
          1958 => x"80", -- $007a6
          1959 => x"7f", -- $007a7
          1960 => x"7f", -- $007a8
          1961 => x"80", -- $007a9
          1962 => x"80", -- $007aa
          1963 => x"80", -- $007ab
          1964 => x"7f", -- $007ac
          1965 => x"7f", -- $007ad
          1966 => x"7f", -- $007ae
          1967 => x"7f", -- $007af
          1968 => x"80", -- $007b0
          1969 => x"80", -- $007b1
          1970 => x"80", -- $007b2
          1971 => x"7f", -- $007b3
          1972 => x"80", -- $007b4
          1973 => x"7f", -- $007b5
          1974 => x"7f", -- $007b6
          1975 => x"7f", -- $007b7
          1976 => x"80", -- $007b8
          1977 => x"80", -- $007b9
          1978 => x"80", -- $007ba
          1979 => x"80", -- $007bb
          1980 => x"80", -- $007bc
          1981 => x"80", -- $007bd
          1982 => x"80", -- $007be
          1983 => x"80", -- $007bf
          1984 => x"80", -- $007c0
          1985 => x"80", -- $007c1
          1986 => x"80", -- $007c2
          1987 => x"80", -- $007c3
          1988 => x"80", -- $007c4
          1989 => x"7f", -- $007c5
          1990 => x"7f", -- $007c6
          1991 => x"7f", -- $007c7
          1992 => x"80", -- $007c8
          1993 => x"80", -- $007c9
          1994 => x"80", -- $007ca
          1995 => x"80", -- $007cb
          1996 => x"80", -- $007cc
          1997 => x"80", -- $007cd
          1998 => x"7f", -- $007ce
          1999 => x"7f", -- $007cf
          2000 => x"7f", -- $007d0
          2001 => x"80", -- $007d1
          2002 => x"80", -- $007d2
          2003 => x"80", -- $007d3
          2004 => x"80", -- $007d4
          2005 => x"7f", -- $007d5
          2006 => x"7f", -- $007d6
          2007 => x"80", -- $007d7
          2008 => x"80", -- $007d8
          2009 => x"80", -- $007d9
          2010 => x"80", -- $007da
          2011 => x"80", -- $007db
          2012 => x"80", -- $007dc
          2013 => x"80", -- $007dd
          2014 => x"80", -- $007de
          2015 => x"80", -- $007df
          2016 => x"80", -- $007e0
          2017 => x"80", -- $007e1
          2018 => x"80", -- $007e2
          2019 => x"80", -- $007e3
          2020 => x"7f", -- $007e4
          2021 => x"80", -- $007e5
          2022 => x"80", -- $007e6
          2023 => x"80", -- $007e7
          2024 => x"7f", -- $007e8
          2025 => x"7f", -- $007e9
          2026 => x"80", -- $007ea
          2027 => x"80", -- $007eb
          2028 => x"80", -- $007ec
          2029 => x"80", -- $007ed
          2030 => x"80", -- $007ee
          2031 => x"80", -- $007ef
          2032 => x"80", -- $007f0
          2033 => x"80", -- $007f1
          2034 => x"80", -- $007f2
          2035 => x"80", -- $007f3
          2036 => x"80", -- $007f4
          2037 => x"80", -- $007f5
          2038 => x"80", -- $007f6
          2039 => x"80", -- $007f7
          2040 => x"80", -- $007f8
          2041 => x"80", -- $007f9
          2042 => x"80", -- $007fa
          2043 => x"80", -- $007fb
          2044 => x"80", -- $007fc
          2045 => x"80", -- $007fd
          2046 => x"80", -- $007fe
          2047 => x"80", -- $007ff
          2048 => x"80", -- $00800
          2049 => x"80", -- $00801
          2050 => x"80", -- $00802
          2051 => x"80", -- $00803
          2052 => x"80", -- $00804
          2053 => x"80", -- $00805
          2054 => x"80", -- $00806
          2055 => x"80", -- $00807
          2056 => x"80", -- $00808
          2057 => x"80", -- $00809
          2058 => x"80", -- $0080a
          2059 => x"80", -- $0080b
          2060 => x"80", -- $0080c
          2061 => x"80", -- $0080d
          2062 => x"80", -- $0080e
          2063 => x"80", -- $0080f
          2064 => x"80", -- $00810
          2065 => x"80", -- $00811
          2066 => x"80", -- $00812
          2067 => x"80", -- $00813
          2068 => x"80", -- $00814
          2069 => x"81", -- $00815
          2070 => x"81", -- $00816
          2071 => x"80", -- $00817
          2072 => x"80", -- $00818
          2073 => x"80", -- $00819
          2074 => x"80", -- $0081a
          2075 => x"81", -- $0081b
          2076 => x"81", -- $0081c
          2077 => x"80", -- $0081d
          2078 => x"80", -- $0081e
          2079 => x"80", -- $0081f
          2080 => x"80", -- $00820
          2081 => x"81", -- $00821
          2082 => x"81", -- $00822
          2083 => x"81", -- $00823
          2084 => x"81", -- $00824
          2085 => x"81", -- $00825
          2086 => x"81", -- $00826
          2087 => x"81", -- $00827
          2088 => x"81", -- $00828
          2089 => x"81", -- $00829
          2090 => x"81", -- $0082a
          2091 => x"81", -- $0082b
          2092 => x"81", -- $0082c
          2093 => x"81", -- $0082d
          2094 => x"81", -- $0082e
          2095 => x"81", -- $0082f
          2096 => x"81", -- $00830
          2097 => x"81", -- $00831
          2098 => x"81", -- $00832
          2099 => x"81", -- $00833
          2100 => x"82", -- $00834
          2101 => x"82", -- $00835
          2102 => x"82", -- $00836
          2103 => x"81", -- $00837
          2104 => x"81", -- $00838
          2105 => x"81", -- $00839
          2106 => x"82", -- $0083a
          2107 => x"82", -- $0083b
          2108 => x"81", -- $0083c
          2109 => x"81", -- $0083d
          2110 => x"81", -- $0083e
          2111 => x"81", -- $0083f
          2112 => x"82", -- $00840
          2113 => x"82", -- $00841
          2114 => x"82", -- $00842
          2115 => x"82", -- $00843
          2116 => x"81", -- $00844
          2117 => x"81", -- $00845
          2118 => x"82", -- $00846
          2119 => x"82", -- $00847
          2120 => x"82", -- $00848
          2121 => x"82", -- $00849
          2122 => x"82", -- $0084a
          2123 => x"82", -- $0084b
          2124 => x"83", -- $0084c
          2125 => x"82", -- $0084d
          2126 => x"82", -- $0084e
          2127 => x"82", -- $0084f
          2128 => x"82", -- $00850
          2129 => x"82", -- $00851
          2130 => x"82", -- $00852
          2131 => x"83", -- $00853
          2132 => x"82", -- $00854
          2133 => x"82", -- $00855
          2134 => x"82", -- $00856
          2135 => x"82", -- $00857
          2136 => x"83", -- $00858
          2137 => x"83", -- $00859
          2138 => x"83", -- $0085a
          2139 => x"83", -- $0085b
          2140 => x"83", -- $0085c
          2141 => x"83", -- $0085d
          2142 => x"83", -- $0085e
          2143 => x"83", -- $0085f
          2144 => x"83", -- $00860
          2145 => x"83", -- $00861
          2146 => x"83", -- $00862
          2147 => x"83", -- $00863
          2148 => x"83", -- $00864
          2149 => x"83", -- $00865
          2150 => x"83", -- $00866
          2151 => x"83", -- $00867
          2152 => x"83", -- $00868
          2153 => x"84", -- $00869
          2154 => x"84", -- $0086a
          2155 => x"84", -- $0086b
          2156 => x"83", -- $0086c
          2157 => x"83", -- $0086d
          2158 => x"84", -- $0086e
          2159 => x"84", -- $0086f
          2160 => x"84", -- $00870
          2161 => x"84", -- $00871
          2162 => x"84", -- $00872
          2163 => x"84", -- $00873
          2164 => x"84", -- $00874
          2165 => x"84", -- $00875
          2166 => x"84", -- $00876
          2167 => x"84", -- $00877
          2168 => x"84", -- $00878
          2169 => x"84", -- $00879
          2170 => x"84", -- $0087a
          2171 => x"85", -- $0087b
          2172 => x"84", -- $0087c
          2173 => x"84", -- $0087d
          2174 => x"84", -- $0087e
          2175 => x"84", -- $0087f
          2176 => x"84", -- $00880
          2177 => x"85", -- $00881
          2178 => x"85", -- $00882
          2179 => x"84", -- $00883
          2180 => x"84", -- $00884
          2181 => x"84", -- $00885
          2182 => x"84", -- $00886
          2183 => x"84", -- $00887
          2184 => x"85", -- $00888
          2185 => x"84", -- $00889
          2186 => x"84", -- $0088a
          2187 => x"84", -- $0088b
          2188 => x"84", -- $0088c
          2189 => x"85", -- $0088d
          2190 => x"85", -- $0088e
          2191 => x"84", -- $0088f
          2192 => x"84", -- $00890
          2193 => x"84", -- $00891
          2194 => x"84", -- $00892
          2195 => x"85", -- $00893
          2196 => x"85", -- $00894
          2197 => x"85", -- $00895
          2198 => x"84", -- $00896
          2199 => x"84", -- $00897
          2200 => x"84", -- $00898
          2201 => x"84", -- $00899
          2202 => x"84", -- $0089a
          2203 => x"84", -- $0089b
          2204 => x"84", -- $0089c
          2205 => x"84", -- $0089d
          2206 => x"84", -- $0089e
          2207 => x"84", -- $0089f
          2208 => x"84", -- $008a0
          2209 => x"84", -- $008a1
          2210 => x"84", -- $008a2
          2211 => x"84", -- $008a3
          2212 => x"84", -- $008a4
          2213 => x"84", -- $008a5
          2214 => x"83", -- $008a6
          2215 => x"84", -- $008a7
          2216 => x"84", -- $008a8
          2217 => x"84", -- $008a9
          2218 => x"84", -- $008aa
          2219 => x"84", -- $008ab
          2220 => x"84", -- $008ac
          2221 => x"83", -- $008ad
          2222 => x"83", -- $008ae
          2223 => x"84", -- $008af
          2224 => x"83", -- $008b0
          2225 => x"83", -- $008b1
          2226 => x"83", -- $008b2
          2227 => x"83", -- $008b3
          2228 => x"84", -- $008b4
          2229 => x"84", -- $008b5
          2230 => x"84", -- $008b6
          2231 => x"84", -- $008b7
          2232 => x"84", -- $008b8
          2233 => x"84", -- $008b9
          2234 => x"84", -- $008ba
          2235 => x"84", -- $008bb
          2236 => x"84", -- $008bc
          2237 => x"84", -- $008bd
          2238 => x"84", -- $008be
          2239 => x"83", -- $008bf
          2240 => x"83", -- $008c0
          2241 => x"84", -- $008c1
          2242 => x"84", -- $008c2
          2243 => x"84", -- $008c3
          2244 => x"84", -- $008c4
          2245 => x"84", -- $008c5
          2246 => x"84", -- $008c6
          2247 => x"83", -- $008c7
          2248 => x"83", -- $008c8
          2249 => x"84", -- $008c9
          2250 => x"84", -- $008ca
          2251 => x"84", -- $008cb
          2252 => x"83", -- $008cc
          2253 => x"83", -- $008cd
          2254 => x"83", -- $008ce
          2255 => x"83", -- $008cf
          2256 => x"83", -- $008d0
          2257 => x"83", -- $008d1
          2258 => x"83", -- $008d2
          2259 => x"83", -- $008d3
          2260 => x"83", -- $008d4
          2261 => x"83", -- $008d5
          2262 => x"83", -- $008d6
          2263 => x"83", -- $008d7
          2264 => x"83", -- $008d8
          2265 => x"83", -- $008d9
          2266 => x"83", -- $008da
          2267 => x"83", -- $008db
          2268 => x"83", -- $008dc
          2269 => x"83", -- $008dd
          2270 => x"83", -- $008de
          2271 => x"83", -- $008df
          2272 => x"83", -- $008e0
          2273 => x"83", -- $008e1
          2274 => x"83", -- $008e2
          2275 => x"83", -- $008e3
          2276 => x"82", -- $008e4
          2277 => x"83", -- $008e5
          2278 => x"83", -- $008e6
          2279 => x"83", -- $008e7
          2280 => x"82", -- $008e8
          2281 => x"82", -- $008e9
          2282 => x"82", -- $008ea
          2283 => x"82", -- $008eb
          2284 => x"83", -- $008ec
          2285 => x"83", -- $008ed
          2286 => x"82", -- $008ee
          2287 => x"82", -- $008ef
          2288 => x"82", -- $008f0
          2289 => x"82", -- $008f1
          2290 => x"82", -- $008f2
          2291 => x"82", -- $008f3
          2292 => x"82", -- $008f4
          2293 => x"82", -- $008f5
          2294 => x"82", -- $008f6
          2295 => x"82", -- $008f7
          2296 => x"82", -- $008f8
          2297 => x"82", -- $008f9
          2298 => x"82", -- $008fa
          2299 => x"82", -- $008fb
          2300 => x"82", -- $008fc
          2301 => x"81", -- $008fd
          2302 => x"81", -- $008fe
          2303 => x"82", -- $008ff
          2304 => x"82", -- $00900
          2305 => x"82", -- $00901
          2306 => x"82", -- $00902
          2307 => x"82", -- $00903
          2308 => x"81", -- $00904
          2309 => x"82", -- $00905
          2310 => x"82", -- $00906
          2311 => x"82", -- $00907
          2312 => x"82", -- $00908
          2313 => x"82", -- $00909
          2314 => x"82", -- $0090a
          2315 => x"82", -- $0090b
          2316 => x"82", -- $0090c
          2317 => x"82", -- $0090d
          2318 => x"82", -- $0090e
          2319 => x"82", -- $0090f
          2320 => x"82", -- $00910
          2321 => x"82", -- $00911
          2322 => x"82", -- $00912
          2323 => x"82", -- $00913
          2324 => x"82", -- $00914
          2325 => x"82", -- $00915
          2326 => x"82", -- $00916
          2327 => x"82", -- $00917
          2328 => x"82", -- $00918
          2329 => x"82", -- $00919
          2330 => x"82", -- $0091a
          2331 => x"82", -- $0091b
          2332 => x"82", -- $0091c
          2333 => x"82", -- $0091d
          2334 => x"82", -- $0091e
          2335 => x"83", -- $0091f
          2336 => x"83", -- $00920
          2337 => x"83", -- $00921
          2338 => x"82", -- $00922
          2339 => x"82", -- $00923
          2340 => x"82", -- $00924
          2341 => x"82", -- $00925
          2342 => x"82", -- $00926
          2343 => x"82", -- $00927
          2344 => x"82", -- $00928
          2345 => x"82", -- $00929
          2346 => x"82", -- $0092a
          2347 => x"83", -- $0092b
          2348 => x"83", -- $0092c
          2349 => x"83", -- $0092d
          2350 => x"82", -- $0092e
          2351 => x"82", -- $0092f
          2352 => x"82", -- $00930
          2353 => x"83", -- $00931
          2354 => x"83", -- $00932
          2355 => x"83", -- $00933
          2356 => x"82", -- $00934
          2357 => x"82", -- $00935
          2358 => x"82", -- $00936
          2359 => x"82", -- $00937
          2360 => x"82", -- $00938
          2361 => x"82", -- $00939
          2362 => x"82", -- $0093a
          2363 => x"82", -- $0093b
          2364 => x"82", -- $0093c
          2365 => x"82", -- $0093d
          2366 => x"82", -- $0093e
          2367 => x"82", -- $0093f
          2368 => x"82", -- $00940
          2369 => x"82", -- $00941
          2370 => x"82", -- $00942
          2371 => x"82", -- $00943
          2372 => x"82", -- $00944
          2373 => x"82", -- $00945
          2374 => x"82", -- $00946
          2375 => x"82", -- $00947
          2376 => x"82", -- $00948
          2377 => x"82", -- $00949
          2378 => x"82", -- $0094a
          2379 => x"81", -- $0094b
          2380 => x"81", -- $0094c
          2381 => x"81", -- $0094d
          2382 => x"81", -- $0094e
          2383 => x"81", -- $0094f
          2384 => x"81", -- $00950
          2385 => x"81", -- $00951
          2386 => x"81", -- $00952
          2387 => x"81", -- $00953
          2388 => x"81", -- $00954
          2389 => x"81", -- $00955
          2390 => x"81", -- $00956
          2391 => x"81", -- $00957
          2392 => x"81", -- $00958
          2393 => x"81", -- $00959
          2394 => x"81", -- $0095a
          2395 => x"81", -- $0095b
          2396 => x"81", -- $0095c
          2397 => x"81", -- $0095d
          2398 => x"81", -- $0095e
          2399 => x"80", -- $0095f
          2400 => x"80", -- $00960
          2401 => x"81", -- $00961
          2402 => x"81", -- $00962
          2403 => x"81", -- $00963
          2404 => x"81", -- $00964
          2405 => x"80", -- $00965
          2406 => x"80", -- $00966
          2407 => x"80", -- $00967
          2408 => x"80", -- $00968
          2409 => x"80", -- $00969
          2410 => x"80", -- $0096a
          2411 => x"80", -- $0096b
          2412 => x"80", -- $0096c
          2413 => x"80", -- $0096d
          2414 => x"80", -- $0096e
          2415 => x"80", -- $0096f
          2416 => x"80", -- $00970
          2417 => x"80", -- $00971
          2418 => x"80", -- $00972
          2419 => x"80", -- $00973
          2420 => x"80", -- $00974
          2421 => x"80", -- $00975
          2422 => x"80", -- $00976
          2423 => x"80", -- $00977
          2424 => x"80", -- $00978
          2425 => x"80", -- $00979
          2426 => x"80", -- $0097a
          2427 => x"80", -- $0097b
          2428 => x"80", -- $0097c
          2429 => x"80", -- $0097d
          2430 => x"80", -- $0097e
          2431 => x"80", -- $0097f
          2432 => x"80", -- $00980
          2433 => x"80", -- $00981
          2434 => x"80", -- $00982
          2435 => x"80", -- $00983
          2436 => x"80", -- $00984
          2437 => x"80", -- $00985
          2438 => x"80", -- $00986
          2439 => x"80", -- $00987
          2440 => x"80", -- $00988
          2441 => x"80", -- $00989
          2442 => x"80", -- $0098a
          2443 => x"80", -- $0098b
          2444 => x"80", -- $0098c
          2445 => x"80", -- $0098d
          2446 => x"80", -- $0098e
          2447 => x"80", -- $0098f
          2448 => x"80", -- $00990
          2449 => x"80", -- $00991
          2450 => x"80", -- $00992
          2451 => x"80", -- $00993
          2452 => x"80", -- $00994
          2453 => x"80", -- $00995
          2454 => x"80", -- $00996
          2455 => x"80", -- $00997
          2456 => x"80", -- $00998
          2457 => x"80", -- $00999
          2458 => x"80", -- $0099a
          2459 => x"80", -- $0099b
          2460 => x"80", -- $0099c
          2461 => x"80", -- $0099d
          2462 => x"7f", -- $0099e
          2463 => x"7f", -- $0099f
          2464 => x"7f", -- $009a0
          2465 => x"7f", -- $009a1
          2466 => x"7f", -- $009a2
          2467 => x"7f", -- $009a3
          2468 => x"7f", -- $009a4
          2469 => x"7f", -- $009a5
          2470 => x"7f", -- $009a6
          2471 => x"7f", -- $009a7
          2472 => x"7f", -- $009a8
          2473 => x"7f", -- $009a9
          2474 => x"7f", -- $009aa
          2475 => x"7f", -- $009ab
          2476 => x"7f", -- $009ac
          2477 => x"7f", -- $009ad
          2478 => x"7f", -- $009ae
          2479 => x"7f", -- $009af
          2480 => x"7f", -- $009b0
          2481 => x"7f", -- $009b1
          2482 => x"7f", -- $009b2
          2483 => x"7e", -- $009b3
          2484 => x"7e", -- $009b4
          2485 => x"7f", -- $009b5
          2486 => x"7f", -- $009b6
          2487 => x"7f", -- $009b7
          2488 => x"7e", -- $009b8
          2489 => x"7e", -- $009b9
          2490 => x"7e", -- $009ba
          2491 => x"7f", -- $009bb
          2492 => x"7f", -- $009bc
          2493 => x"7f", -- $009bd
          2494 => x"7f", -- $009be
          2495 => x"7e", -- $009bf
          2496 => x"7e", -- $009c0
          2497 => x"7e", -- $009c1
          2498 => x"7e", -- $009c2
          2499 => x"7e", -- $009c3
          2500 => x"7e", -- $009c4
          2501 => x"7e", -- $009c5
          2502 => x"7e", -- $009c6
          2503 => x"7e", -- $009c7
          2504 => x"7e", -- $009c8
          2505 => x"7e", -- $009c9
          2506 => x"7e", -- $009ca
          2507 => x"7e", -- $009cb
          2508 => x"7e", -- $009cc
          2509 => x"7e", -- $009cd
          2510 => x"7e", -- $009ce
          2511 => x"7e", -- $009cf
          2512 => x"7e", -- $009d0
          2513 => x"7e", -- $009d1
          2514 => x"7e", -- $009d2
          2515 => x"7e", -- $009d3
          2516 => x"7e", -- $009d4
          2517 => x"7e", -- $009d5
          2518 => x"7e", -- $009d6
          2519 => x"7e", -- $009d7
          2520 => x"7e", -- $009d8
          2521 => x"7e", -- $009d9
          2522 => x"7e", -- $009da
          2523 => x"7e", -- $009db
          2524 => x"7e", -- $009dc
          2525 => x"7e", -- $009dd
          2526 => x"7e", -- $009de
          2527 => x"7e", -- $009df
          2528 => x"7e", -- $009e0
          2529 => x"7e", -- $009e1
          2530 => x"7e", -- $009e2
          2531 => x"7e", -- $009e3
          2532 => x"7e", -- $009e4
          2533 => x"7e", -- $009e5
          2534 => x"7e", -- $009e6
          2535 => x"7e", -- $009e7
          2536 => x"7e", -- $009e8
          2537 => x"7e", -- $009e9
          2538 => x"7e", -- $009ea
          2539 => x"7e", -- $009eb
          2540 => x"7e", -- $009ec
          2541 => x"7e", -- $009ed
          2542 => x"7e", -- $009ee
          2543 => x"7e", -- $009ef
          2544 => x"7e", -- $009f0
          2545 => x"7e", -- $009f1
          2546 => x"7e", -- $009f2
          2547 => x"7e", -- $009f3
          2548 => x"7e", -- $009f4
          2549 => x"7e", -- $009f5
          2550 => x"7e", -- $009f6
          2551 => x"7e", -- $009f7
          2552 => x"7e", -- $009f8
          2553 => x"7e", -- $009f9
          2554 => x"7e", -- $009fa
          2555 => x"7e", -- $009fb
          2556 => x"7e", -- $009fc
          2557 => x"7e", -- $009fd
          2558 => x"7e", -- $009fe
          2559 => x"7e", -- $009ff
          2560 => x"7e", -- $00a00
          2561 => x"7e", -- $00a01
          2562 => x"7e", -- $00a02
          2563 => x"7e", -- $00a03
          2564 => x"7e", -- $00a04
          2565 => x"7e", -- $00a05
          2566 => x"7e", -- $00a06
          2567 => x"7e", -- $00a07
          2568 => x"7e", -- $00a08
          2569 => x"7e", -- $00a09
          2570 => x"7d", -- $00a0a
          2571 => x"7d", -- $00a0b
          2572 => x"7d", -- $00a0c
          2573 => x"7d", -- $00a0d
          2574 => x"7d", -- $00a0e
          2575 => x"7d", -- $00a0f
          2576 => x"7d", -- $00a10
          2577 => x"7d", -- $00a11
          2578 => x"7d", -- $00a12
          2579 => x"7d", -- $00a13
          2580 => x"7d", -- $00a14
          2581 => x"7d", -- $00a15
          2582 => x"7d", -- $00a16
          2583 => x"7d", -- $00a17
          2584 => x"7d", -- $00a18
          2585 => x"7d", -- $00a19
          2586 => x"7d", -- $00a1a
          2587 => x"7d", -- $00a1b
          2588 => x"7d", -- $00a1c
          2589 => x"7d", -- $00a1d
          2590 => x"7d", -- $00a1e
          2591 => x"7d", -- $00a1f
          2592 => x"7d", -- $00a20
          2593 => x"7d", -- $00a21
          2594 => x"7d", -- $00a22
          2595 => x"7d", -- $00a23
          2596 => x"7d", -- $00a24
          2597 => x"7d", -- $00a25
          2598 => x"7d", -- $00a26
          2599 => x"7d", -- $00a27
          2600 => x"7d", -- $00a28
          2601 => x"7d", -- $00a29
          2602 => x"7d", -- $00a2a
          2603 => x"7d", -- $00a2b
          2604 => x"7d", -- $00a2c
          2605 => x"7d", -- $00a2d
          2606 => x"7d", -- $00a2e
          2607 => x"7c", -- $00a2f
          2608 => x"7d", -- $00a30
          2609 => x"7d", -- $00a31
          2610 => x"7d", -- $00a32
          2611 => x"7d", -- $00a33
          2612 => x"7d", -- $00a34
          2613 => x"7c", -- $00a35
          2614 => x"7d", -- $00a36
          2615 => x"7c", -- $00a37
          2616 => x"7c", -- $00a38
          2617 => x"7c", -- $00a39
          2618 => x"7d", -- $00a3a
          2619 => x"7d", -- $00a3b
          2620 => x"7c", -- $00a3c
          2621 => x"7c", -- $00a3d
          2622 => x"7c", -- $00a3e
          2623 => x"7c", -- $00a3f
          2624 => x"7c", -- $00a40
          2625 => x"7c", -- $00a41
          2626 => x"7c", -- $00a42
          2627 => x"7c", -- $00a43
          2628 => x"7c", -- $00a44
          2629 => x"7c", -- $00a45
          2630 => x"7c", -- $00a46
          2631 => x"7c", -- $00a47
          2632 => x"7c", -- $00a48
          2633 => x"7c", -- $00a49
          2634 => x"7d", -- $00a4a
          2635 => x"7d", -- $00a4b
          2636 => x"7d", -- $00a4c
          2637 => x"7d", -- $00a4d
          2638 => x"7d", -- $00a4e
          2639 => x"7d", -- $00a4f
          2640 => x"7d", -- $00a50
          2641 => x"7c", -- $00a51
          2642 => x"7c", -- $00a52
          2643 => x"7c", -- $00a53
          2644 => x"7d", -- $00a54
          2645 => x"7d", -- $00a55
          2646 => x"7d", -- $00a56
          2647 => x"7d", -- $00a57
          2648 => x"7d", -- $00a58
          2649 => x"7d", -- $00a59
          2650 => x"7d", -- $00a5a
          2651 => x"7d", -- $00a5b
          2652 => x"7d", -- $00a5c
          2653 => x"7d", -- $00a5d
          2654 => x"7d", -- $00a5e
          2655 => x"7d", -- $00a5f
          2656 => x"7d", -- $00a60
          2657 => x"7d", -- $00a61
          2658 => x"7d", -- $00a62
          2659 => x"7d", -- $00a63
          2660 => x"7d", -- $00a64
          2661 => x"7d", -- $00a65
          2662 => x"7d", -- $00a66
          2663 => x"7d", -- $00a67
          2664 => x"7d", -- $00a68
          2665 => x"7d", -- $00a69
          2666 => x"7d", -- $00a6a
          2667 => x"7d", -- $00a6b
          2668 => x"7d", -- $00a6c
          2669 => x"7d", -- $00a6d
          2670 => x"7d", -- $00a6e
          2671 => x"7d", -- $00a6f
          2672 => x"7d", -- $00a70
          2673 => x"7d", -- $00a71
          2674 => x"7d", -- $00a72
          2675 => x"7d", -- $00a73
          2676 => x"7d", -- $00a74
          2677 => x"7d", -- $00a75
          2678 => x"7d", -- $00a76
          2679 => x"7d", -- $00a77
          2680 => x"7d", -- $00a78
          2681 => x"7d", -- $00a79
          2682 => x"7d", -- $00a7a
          2683 => x"7d", -- $00a7b
          2684 => x"7d", -- $00a7c
          2685 => x"7d", -- $00a7d
          2686 => x"7d", -- $00a7e
          2687 => x"7d", -- $00a7f
          2688 => x"7d", -- $00a80
          2689 => x"7d", -- $00a81
          2690 => x"7d", -- $00a82
          2691 => x"7d", -- $00a83
          2692 => x"7d", -- $00a84
          2693 => x"7d", -- $00a85
          2694 => x"7d", -- $00a86
          2695 => x"7d", -- $00a87
          2696 => x"7d", -- $00a88
          2697 => x"7d", -- $00a89
          2698 => x"7e", -- $00a8a
          2699 => x"7d", -- $00a8b
          2700 => x"7d", -- $00a8c
          2701 => x"7e", -- $00a8d
          2702 => x"7e", -- $00a8e
          2703 => x"7e", -- $00a8f
          2704 => x"7d", -- $00a90
          2705 => x"7d", -- $00a91
          2706 => x"7d", -- $00a92
          2707 => x"7d", -- $00a93
          2708 => x"7e", -- $00a94
          2709 => x"7e", -- $00a95
          2710 => x"7e", -- $00a96
          2711 => x"7e", -- $00a97
          2712 => x"7e", -- $00a98
          2713 => x"7e", -- $00a99
          2714 => x"7e", -- $00a9a
          2715 => x"7e", -- $00a9b
          2716 => x"7e", -- $00a9c
          2717 => x"7e", -- $00a9d
          2718 => x"7e", -- $00a9e
          2719 => x"7e", -- $00a9f
          2720 => x"7e", -- $00aa0
          2721 => x"7e", -- $00aa1
          2722 => x"7e", -- $00aa2
          2723 => x"7e", -- $00aa3
          2724 => x"7e", -- $00aa4
          2725 => x"7e", -- $00aa5
          2726 => x"7e", -- $00aa6
          2727 => x"7e", -- $00aa7
          2728 => x"7e", -- $00aa8
          2729 => x"7e", -- $00aa9
          2730 => x"7e", -- $00aaa
          2731 => x"7e", -- $00aab
          2732 => x"7e", -- $00aac
          2733 => x"7e", -- $00aad
          2734 => x"7e", -- $00aae
          2735 => x"7e", -- $00aaf
          2736 => x"7e", -- $00ab0
          2737 => x"7f", -- $00ab1
          2738 => x"7f", -- $00ab2
          2739 => x"7f", -- $00ab3
          2740 => x"7f", -- $00ab4
          2741 => x"7f", -- $00ab5
          2742 => x"7f", -- $00ab6
          2743 => x"7f", -- $00ab7
          2744 => x"7e", -- $00ab8
          2745 => x"7f", -- $00ab9
          2746 => x"7f", -- $00aba
          2747 => x"7f", -- $00abb
          2748 => x"7f", -- $00abc
          2749 => x"7f", -- $00abd
          2750 => x"7f", -- $00abe
          2751 => x"7f", -- $00abf
          2752 => x"7f", -- $00ac0
          2753 => x"7f", -- $00ac1
          2754 => x"7f", -- $00ac2
          2755 => x"7f", -- $00ac3
          2756 => x"7f", -- $00ac4
          2757 => x"7f", -- $00ac5
          2758 => x"7f", -- $00ac6
          2759 => x"7f", -- $00ac7
          2760 => x"7f", -- $00ac8
          2761 => x"7f", -- $00ac9
          2762 => x"7f", -- $00aca
          2763 => x"7f", -- $00acb
          2764 => x"7f", -- $00acc
          2765 => x"7f", -- $00acd
          2766 => x"7f", -- $00ace
          2767 => x"7f", -- $00acf
          2768 => x"7f", -- $00ad0
          2769 => x"7f", -- $00ad1
          2770 => x"7f", -- $00ad2
          2771 => x"7f", -- $00ad3
          2772 => x"7f", -- $00ad4
          2773 => x"7f", -- $00ad5
          2774 => x"7f", -- $00ad6
          2775 => x"7f", -- $00ad7
          2776 => x"7f", -- $00ad8
          2777 => x"7f", -- $00ad9
          2778 => x"80", -- $00ada
          2779 => x"80", -- $00adb
          2780 => x"7f", -- $00adc
          2781 => x"7f", -- $00add
          2782 => x"80", -- $00ade
          2783 => x"80", -- $00adf
          2784 => x"7f", -- $00ae0
          2785 => x"7f", -- $00ae1
          2786 => x"7f", -- $00ae2
          2787 => x"80", -- $00ae3
          2788 => x"80", -- $00ae4
          2789 => x"80", -- $00ae5
          2790 => x"80", -- $00ae6
          2791 => x"80", -- $00ae7
          2792 => x"80", -- $00ae8
          2793 => x"80", -- $00ae9
          2794 => x"80", -- $00aea
          2795 => x"80", -- $00aeb
          2796 => x"80", -- $00aec
          2797 => x"80", -- $00aed
          2798 => x"80", -- $00aee
          2799 => x"80", -- $00aef
          2800 => x"80", -- $00af0
          2801 => x"80", -- $00af1
          2802 => x"80", -- $00af2
          2803 => x"80", -- $00af3
          2804 => x"80", -- $00af4
          2805 => x"80", -- $00af5
          2806 => x"80", -- $00af6
          2807 => x"80", -- $00af7
          2808 => x"80", -- $00af8
          2809 => x"80", -- $00af9
          2810 => x"80", -- $00afa
          2811 => x"80", -- $00afb
          2812 => x"80", -- $00afc
          2813 => x"80", -- $00afd
          2814 => x"80", -- $00afe
          2815 => x"80", -- $00aff
          2816 => x"80", -- $00b00
          2817 => x"80", -- $00b01
          2818 => x"80", -- $00b02
          2819 => x"80", -- $00b03
          2820 => x"80", -- $00b04
          2821 => x"80", -- $00b05
          2822 => x"80", -- $00b06
          2823 => x"80", -- $00b07
          2824 => x"80", -- $00b08
          2825 => x"80", -- $00b09
          2826 => x"80", -- $00b0a
          2827 => x"80", -- $00b0b
          2828 => x"80", -- $00b0c
          2829 => x"80", -- $00b0d
          2830 => x"80", -- $00b0e
          2831 => x"80", -- $00b0f
          2832 => x"80", -- $00b10
          2833 => x"80", -- $00b11
          2834 => x"80", -- $00b12
          2835 => x"80", -- $00b13
          2836 => x"80", -- $00b14
          2837 => x"81", -- $00b15
          2838 => x"81", -- $00b16
          2839 => x"81", -- $00b17
          2840 => x"81", -- $00b18
          2841 => x"81", -- $00b19
          2842 => x"81", -- $00b1a
          2843 => x"81", -- $00b1b
          2844 => x"81", -- $00b1c
          2845 => x"81", -- $00b1d
          2846 => x"81", -- $00b1e
          2847 => x"81", -- $00b1f
          2848 => x"81", -- $00b20
          2849 => x"81", -- $00b21
          2850 => x"81", -- $00b22
          2851 => x"81", -- $00b23
          2852 => x"81", -- $00b24
          2853 => x"81", -- $00b25
          2854 => x"81", -- $00b26
          2855 => x"81", -- $00b27
          2856 => x"81", -- $00b28
          2857 => x"81", -- $00b29
          2858 => x"82", -- $00b2a
          2859 => x"82", -- $00b2b
          2860 => x"82", -- $00b2c
          2861 => x"82", -- $00b2d
          2862 => x"82", -- $00b2e
          2863 => x"82", -- $00b2f
          2864 => x"82", -- $00b30
          2865 => x"82", -- $00b31
          2866 => x"82", -- $00b32
          2867 => x"82", -- $00b33
          2868 => x"82", -- $00b34
          2869 => x"82", -- $00b35
          2870 => x"82", -- $00b36
          2871 => x"82", -- $00b37
          2872 => x"82", -- $00b38
          2873 => x"82", -- $00b39
          2874 => x"82", -- $00b3a
          2875 => x"82", -- $00b3b
          2876 => x"82", -- $00b3c
          2877 => x"82", -- $00b3d
          2878 => x"82", -- $00b3e
          2879 => x"82", -- $00b3f
          2880 => x"82", -- $00b40
          2881 => x"82", -- $00b41
          2882 => x"82", -- $00b42
          2883 => x"82", -- $00b43
          2884 => x"82", -- $00b44
          2885 => x"82", -- $00b45
          2886 => x"82", -- $00b46
          2887 => x"82", -- $00b47
          2888 => x"82", -- $00b48
          2889 => x"82", -- $00b49
          2890 => x"82", -- $00b4a
          2891 => x"82", -- $00b4b
          2892 => x"82", -- $00b4c
          2893 => x"82", -- $00b4d
          2894 => x"82", -- $00b4e
          2895 => x"82", -- $00b4f
          2896 => x"82", -- $00b50
          2897 => x"82", -- $00b51
          2898 => x"82", -- $00b52
          2899 => x"82", -- $00b53
          2900 => x"82", -- $00b54
          2901 => x"82", -- $00b55
          2902 => x"82", -- $00b56
          2903 => x"82", -- $00b57
          2904 => x"82", -- $00b58
          2905 => x"82", -- $00b59
          2906 => x"83", -- $00b5a
          2907 => x"82", -- $00b5b
          2908 => x"82", -- $00b5c
          2909 => x"83", -- $00b5d
          2910 => x"83", -- $00b5e
          2911 => x"83", -- $00b5f
          2912 => x"83", -- $00b60
          2913 => x"83", -- $00b61
          2914 => x"83", -- $00b62
          2915 => x"82", -- $00b63
          2916 => x"83", -- $00b64
          2917 => x"83", -- $00b65
          2918 => x"83", -- $00b66
          2919 => x"83", -- $00b67
          2920 => x"83", -- $00b68
          2921 => x"83", -- $00b69
          2922 => x"83", -- $00b6a
          2923 => x"83", -- $00b6b
          2924 => x"83", -- $00b6c
          2925 => x"83", -- $00b6d
          2926 => x"83", -- $00b6e
          2927 => x"83", -- $00b6f
          2928 => x"83", -- $00b70
          2929 => x"83", -- $00b71
          2930 => x"83", -- $00b72
          2931 => x"83", -- $00b73
          2932 => x"83", -- $00b74
          2933 => x"83", -- $00b75
          2934 => x"83", -- $00b76
          2935 => x"83", -- $00b77
          2936 => x"83", -- $00b78
          2937 => x"83", -- $00b79
          2938 => x"83", -- $00b7a
          2939 => x"83", -- $00b7b
          2940 => x"83", -- $00b7c
          2941 => x"83", -- $00b7d
          2942 => x"83", -- $00b7e
          2943 => x"83", -- $00b7f
          2944 => x"83", -- $00b80
          2945 => x"83", -- $00b81
          2946 => x"83", -- $00b82
          2947 => x"83", -- $00b83
          2948 => x"83", -- $00b84
          2949 => x"83", -- $00b85
          2950 => x"83", -- $00b86
          2951 => x"83", -- $00b87
          2952 => x"83", -- $00b88
          2953 => x"83", -- $00b89
          2954 => x"83", -- $00b8a
          2955 => x"83", -- $00b8b
          2956 => x"83", -- $00b8c
          2957 => x"83", -- $00b8d
          2958 => x"83", -- $00b8e
          2959 => x"83", -- $00b8f
          2960 => x"83", -- $00b90
          2961 => x"83", -- $00b91
          2962 => x"84", -- $00b92
          2963 => x"84", -- $00b93
          2964 => x"84", -- $00b94
          2965 => x"84", -- $00b95
          2966 => x"84", -- $00b96
          2967 => x"84", -- $00b97
          2968 => x"84", -- $00b98
          2969 => x"84", -- $00b99
          2970 => x"84", -- $00b9a
          2971 => x"84", -- $00b9b
          2972 => x"84", -- $00b9c
          2973 => x"84", -- $00b9d
          2974 => x"84", -- $00b9e
          2975 => x"84", -- $00b9f
          2976 => x"84", -- $00ba0
          2977 => x"84", -- $00ba1
          2978 => x"84", -- $00ba2
          2979 => x"84", -- $00ba3
          2980 => x"84", -- $00ba4
          2981 => x"84", -- $00ba5
          2982 => x"84", -- $00ba6
          2983 => x"84", -- $00ba7
          2984 => x"84", -- $00ba8
          2985 => x"84", -- $00ba9
          2986 => x"84", -- $00baa
          2987 => x"84", -- $00bab
          2988 => x"84", -- $00bac
          2989 => x"84", -- $00bad
          2990 => x"84", -- $00bae
          2991 => x"84", -- $00baf
          2992 => x"84", -- $00bb0
          2993 => x"84", -- $00bb1
          2994 => x"84", -- $00bb2
          2995 => x"84", -- $00bb3
          2996 => x"84", -- $00bb4
          2997 => x"84", -- $00bb5
          2998 => x"84", -- $00bb6
          2999 => x"84", -- $00bb7
          3000 => x"84", -- $00bb8
          3001 => x"84", -- $00bb9
          3002 => x"85", -- $00bba
          3003 => x"85", -- $00bbb
          3004 => x"85", -- $00bbc
          3005 => x"84", -- $00bbd
          3006 => x"84", -- $00bbe
          3007 => x"84", -- $00bbf
          3008 => x"84", -- $00bc0
          3009 => x"85", -- $00bc1
          3010 => x"85", -- $00bc2
          3011 => x"85", -- $00bc3
          3012 => x"85", -- $00bc4
          3013 => x"84", -- $00bc5
          3014 => x"84", -- $00bc6
          3015 => x"85", -- $00bc7
          3016 => x"85", -- $00bc8
          3017 => x"85", -- $00bc9
          3018 => x"84", -- $00bca
          3019 => x"84", -- $00bcb
          3020 => x"84", -- $00bcc
          3021 => x"84", -- $00bcd
          3022 => x"84", -- $00bce
          3023 => x"84", -- $00bcf
          3024 => x"85", -- $00bd0
          3025 => x"85", -- $00bd1
          3026 => x"85", -- $00bd2
          3027 => x"85", -- $00bd3
          3028 => x"84", -- $00bd4
          3029 => x"84", -- $00bd5
          3030 => x"84", -- $00bd6
          3031 => x"84", -- $00bd7
          3032 => x"84", -- $00bd8
          3033 => x"84", -- $00bd9
          3034 => x"84", -- $00bda
          3035 => x"84", -- $00bdb
          3036 => x"84", -- $00bdc
          3037 => x"84", -- $00bdd
          3038 => x"84", -- $00bde
          3039 => x"84", -- $00bdf
          3040 => x"84", -- $00be0
          3041 => x"84", -- $00be1
          3042 => x"84", -- $00be2
          3043 => x"84", -- $00be3
          3044 => x"84", -- $00be4
          3045 => x"84", -- $00be5
          3046 => x"84", -- $00be6
          3047 => x"84", -- $00be7
          3048 => x"84", -- $00be8
          3049 => x"84", -- $00be9
          3050 => x"84", -- $00bea
          3051 => x"84", -- $00beb
          3052 => x"84", -- $00bec
          3053 => x"84", -- $00bed
          3054 => x"84", -- $00bee
          3055 => x"84", -- $00bef
          3056 => x"84", -- $00bf0
          3057 => x"84", -- $00bf1
          3058 => x"84", -- $00bf2
          3059 => x"84", -- $00bf3
          3060 => x"84", -- $00bf4
          3061 => x"84", -- $00bf5
          3062 => x"84", -- $00bf6
          3063 => x"84", -- $00bf7
          3064 => x"84", -- $00bf8
          3065 => x"84", -- $00bf9
          3066 => x"84", -- $00bfa
          3067 => x"83", -- $00bfb
          3068 => x"83", -- $00bfc
          3069 => x"83", -- $00bfd
          3070 => x"83", -- $00bfe
          3071 => x"83", -- $00bff
          3072 => x"83", -- $00c00
          3073 => x"83", -- $00c01
          3074 => x"83", -- $00c02
          3075 => x"83", -- $00c03
          3076 => x"83", -- $00c04
          3077 => x"83", -- $00c05
          3078 => x"83", -- $00c06
          3079 => x"83", -- $00c07
          3080 => x"83", -- $00c08
          3081 => x"83", -- $00c09
          3082 => x"83", -- $00c0a
          3083 => x"83", -- $00c0b
          3084 => x"83", -- $00c0c
          3085 => x"83", -- $00c0d
          3086 => x"83", -- $00c0e
          3087 => x"83", -- $00c0f
          3088 => x"83", -- $00c10
          3089 => x"83", -- $00c11
          3090 => x"82", -- $00c12
          3091 => x"82", -- $00c13
          3092 => x"82", -- $00c14
          3093 => x"82", -- $00c15
          3094 => x"82", -- $00c16
          3095 => x"82", -- $00c17
          3096 => x"82", -- $00c18
          3097 => x"82", -- $00c19
          3098 => x"82", -- $00c1a
          3099 => x"82", -- $00c1b
          3100 => x"82", -- $00c1c
          3101 => x"82", -- $00c1d
          3102 => x"82", -- $00c1e
          3103 => x"82", -- $00c1f
          3104 => x"82", -- $00c20
          3105 => x"82", -- $00c21
          3106 => x"82", -- $00c22
          3107 => x"82", -- $00c23
          3108 => x"82", -- $00c24
          3109 => x"82", -- $00c25
          3110 => x"82", -- $00c26
          3111 => x"82", -- $00c27
          3112 => x"82", -- $00c28
          3113 => x"81", -- $00c29
          3114 => x"81", -- $00c2a
          3115 => x"81", -- $00c2b
          3116 => x"81", -- $00c2c
          3117 => x"81", -- $00c2d
          3118 => x"81", -- $00c2e
          3119 => x"81", -- $00c2f
          3120 => x"81", -- $00c30
          3121 => x"81", -- $00c31
          3122 => x"81", -- $00c32
          3123 => x"81", -- $00c33
          3124 => x"81", -- $00c34
          3125 => x"81", -- $00c35
          3126 => x"81", -- $00c36
          3127 => x"81", -- $00c37
          3128 => x"81", -- $00c38
          3129 => x"81", -- $00c39
          3130 => x"81", -- $00c3a
          3131 => x"81", -- $00c3b
          3132 => x"81", -- $00c3c
          3133 => x"81", -- $00c3d
          3134 => x"81", -- $00c3e
          3135 => x"81", -- $00c3f
          3136 => x"80", -- $00c40
          3137 => x"80", -- $00c41
          3138 => x"80", -- $00c42
          3139 => x"80", -- $00c43
          3140 => x"80", -- $00c44
          3141 => x"80", -- $00c45
          3142 => x"80", -- $00c46
          3143 => x"80", -- $00c47
          3144 => x"80", -- $00c48
          3145 => x"80", -- $00c49
          3146 => x"80", -- $00c4a
          3147 => x"80", -- $00c4b
          3148 => x"80", -- $00c4c
          3149 => x"80", -- $00c4d
          3150 => x"80", -- $00c4e
          3151 => x"80", -- $00c4f
          3152 => x"80", -- $00c50
          3153 => x"80", -- $00c51
          3154 => x"80", -- $00c52
          3155 => x"80", -- $00c53
          3156 => x"80", -- $00c54
          3157 => x"80", -- $00c55
          3158 => x"80", -- $00c56
          3159 => x"80", -- $00c57
          3160 => x"80", -- $00c58
          3161 => x"80", -- $00c59
          3162 => x"80", -- $00c5a
          3163 => x"80", -- $00c5b
          3164 => x"80", -- $00c5c
          3165 => x"80", -- $00c5d
          3166 => x"80", -- $00c5e
          3167 => x"80", -- $00c5f
          3168 => x"80", -- $00c60
          3169 => x"80", -- $00c61
          3170 => x"80", -- $00c62
          3171 => x"80", -- $00c63
          3172 => x"80", -- $00c64
          3173 => x"80", -- $00c65
          3174 => x"80", -- $00c66
          3175 => x"80", -- $00c67
          3176 => x"80", -- $00c68
          3177 => x"80", -- $00c69
          3178 => x"80", -- $00c6a
          3179 => x"80", -- $00c6b
          3180 => x"80", -- $00c6c
          3181 => x"80", -- $00c6d
          3182 => x"80", -- $00c6e
          3183 => x"80", -- $00c6f
          3184 => x"80", -- $00c70
          3185 => x"80", -- $00c71
          3186 => x"80", -- $00c72
          3187 => x"80", -- $00c73
          3188 => x"80", -- $00c74
          3189 => x"80", -- $00c75
          3190 => x"80", -- $00c76
          3191 => x"80", -- $00c77
          3192 => x"80", -- $00c78
          3193 => x"80", -- $00c79
          3194 => x"80", -- $00c7a
          3195 => x"80", -- $00c7b
          3196 => x"80", -- $00c7c
          3197 => x"80", -- $00c7d
          3198 => x"80", -- $00c7e
          3199 => x"80", -- $00c7f
          3200 => x"80", -- $00c80
          3201 => x"80", -- $00c81
          3202 => x"80", -- $00c82
          3203 => x"80", -- $00c83
          3204 => x"80", -- $00c84
          3205 => x"80", -- $00c85
          3206 => x"80", -- $00c86
          3207 => x"80", -- $00c87
          3208 => x"80", -- $00c88
          3209 => x"80", -- $00c89
          3210 => x"80", -- $00c8a
          3211 => x"80", -- $00c8b
          3212 => x"80", -- $00c8c
          3213 => x"80", -- $00c8d
          3214 => x"80", -- $00c8e
          3215 => x"80", -- $00c8f
          3216 => x"80", -- $00c90
          3217 => x"80", -- $00c91
          3218 => x"80", -- $00c92
          3219 => x"80", -- $00c93
          3220 => x"80", -- $00c94
          3221 => x"80", -- $00c95
          3222 => x"80", -- $00c96
          3223 => x"80", -- $00c97
          3224 => x"80", -- $00c98
          3225 => x"80", -- $00c99
          3226 => x"80", -- $00c9a
          3227 => x"80", -- $00c9b
          3228 => x"80", -- $00c9c
          3229 => x"80", -- $00c9d
          3230 => x"7f", -- $00c9e
          3231 => x"7f", -- $00c9f
          3232 => x"7f", -- $00ca0
          3233 => x"7f", -- $00ca1
          3234 => x"7f", -- $00ca2
          3235 => x"7f", -- $00ca3
          3236 => x"7f", -- $00ca4
          3237 => x"7f", -- $00ca5
          3238 => x"7f", -- $00ca6
          3239 => x"7f", -- $00ca7
          3240 => x"7f", -- $00ca8
          3241 => x"7f", -- $00ca9
          3242 => x"7f", -- $00caa
          3243 => x"7f", -- $00cab
          3244 => x"7f", -- $00cac
          3245 => x"7f", -- $00cad
          3246 => x"7f", -- $00cae
          3247 => x"7f", -- $00caf
          3248 => x"7f", -- $00cb0
          3249 => x"7f", -- $00cb1
          3250 => x"7f", -- $00cb2
          3251 => x"7f", -- $00cb3
          3252 => x"7f", -- $00cb4
          3253 => x"7f", -- $00cb5
          3254 => x"7f", -- $00cb6
          3255 => x"7f", -- $00cb7
          3256 => x"7f", -- $00cb8
          3257 => x"7f", -- $00cb9
          3258 => x"7f", -- $00cba
          3259 => x"7f", -- $00cbb
          3260 => x"7f", -- $00cbc
          3261 => x"7f", -- $00cbd
          3262 => x"7f", -- $00cbe
          3263 => x"7f", -- $00cbf
          3264 => x"7e", -- $00cc0
          3265 => x"7f", -- $00cc1
          3266 => x"7e", -- $00cc2
          3267 => x"7e", -- $00cc3
          3268 => x"7e", -- $00cc4
          3269 => x"7e", -- $00cc5
          3270 => x"7e", -- $00cc6
          3271 => x"7e", -- $00cc7
          3272 => x"7e", -- $00cc8
          3273 => x"7e", -- $00cc9
          3274 => x"7e", -- $00cca
          3275 => x"7e", -- $00ccb
          3276 => x"7e", -- $00ccc
          3277 => x"7e", -- $00ccd
          3278 => x"7e", -- $00cce
          3279 => x"7e", -- $00ccf
          3280 => x"7e", -- $00cd0
          3281 => x"7e", -- $00cd1
          3282 => x"7e", -- $00cd2
          3283 => x"7e", -- $00cd3
          3284 => x"7e", -- $00cd4
          3285 => x"7e", -- $00cd5
          3286 => x"7e", -- $00cd6
          3287 => x"7e", -- $00cd7
          3288 => x"7e", -- $00cd8
          3289 => x"7e", -- $00cd9
          3290 => x"7e", -- $00cda
          3291 => x"7e", -- $00cdb
          3292 => x"7e", -- $00cdc
          3293 => x"7e", -- $00cdd
          3294 => x"7e", -- $00cde
          3295 => x"7e", -- $00cdf
          3296 => x"7e", -- $00ce0
          3297 => x"7e", -- $00ce1
          3298 => x"7e", -- $00ce2
          3299 => x"7e", -- $00ce3
          3300 => x"7e", -- $00ce4
          3301 => x"7e", -- $00ce5
          3302 => x"7e", -- $00ce6
          3303 => x"7e", -- $00ce7
          3304 => x"7e", -- $00ce8
          3305 => x"7e", -- $00ce9
          3306 => x"7e", -- $00cea
          3307 => x"7e", -- $00ceb
          3308 => x"7e", -- $00cec
          3309 => x"7e", -- $00ced
          3310 => x"7d", -- $00cee
          3311 => x"7d", -- $00cef
          3312 => x"7e", -- $00cf0
          3313 => x"7e", -- $00cf1
          3314 => x"7e", -- $00cf2
          3315 => x"7e", -- $00cf3
          3316 => x"7e", -- $00cf4
          3317 => x"7e", -- $00cf5
          3318 => x"7d", -- $00cf6
          3319 => x"7e", -- $00cf7
          3320 => x"7e", -- $00cf8
          3321 => x"7e", -- $00cf9
          3322 => x"7d", -- $00cfa
          3323 => x"7d", -- $00cfb
          3324 => x"7d", -- $00cfc
          3325 => x"7d", -- $00cfd
          3326 => x"7d", -- $00cfe
          3327 => x"7d", -- $00cff
          3328 => x"7d", -- $00d00
          3329 => x"7e", -- $00d01
          3330 => x"7d", -- $00d02
          3331 => x"7d", -- $00d03
          3332 => x"7d", -- $00d04
          3333 => x"7d", -- $00d05
          3334 => x"7d", -- $00d06
          3335 => x"7d", -- $00d07
          3336 => x"7d", -- $00d08
          3337 => x"7d", -- $00d09
          3338 => x"7d", -- $00d0a
          3339 => x"7d", -- $00d0b
          3340 => x"7d", -- $00d0c
          3341 => x"7d", -- $00d0d
          3342 => x"7d", -- $00d0e
          3343 => x"7d", -- $00d0f
          3344 => x"7d", -- $00d10
          3345 => x"7d", -- $00d11
          3346 => x"7d", -- $00d12
          3347 => x"7c", -- $00d13
          3348 => x"7d", -- $00d14
          3349 => x"7d", -- $00d15
          3350 => x"7d", -- $00d16
          3351 => x"7d", -- $00d17
          3352 => x"7d", -- $00d18
          3353 => x"7d", -- $00d19
          3354 => x"7d", -- $00d1a
          3355 => x"7d", -- $00d1b
          3356 => x"7c", -- $00d1c
          3357 => x"7c", -- $00d1d
          3358 => x"7c", -- $00d1e
          3359 => x"7c", -- $00d1f
          3360 => x"7c", -- $00d20
          3361 => x"7c", -- $00d21
          3362 => x"7c", -- $00d22
          3363 => x"7c", -- $00d23
          3364 => x"7c", -- $00d24
          3365 => x"7c", -- $00d25
          3366 => x"7d", -- $00d26
          3367 => x"7d", -- $00d27
          3368 => x"7d", -- $00d28
          3369 => x"7d", -- $00d29
          3370 => x"7d", -- $00d2a
          3371 => x"7c", -- $00d2b
          3372 => x"7c", -- $00d2c
          3373 => x"7c", -- $00d2d
          3374 => x"7c", -- $00d2e
          3375 => x"7c", -- $00d2f
          3376 => x"7d", -- $00d30
          3377 => x"7d", -- $00d31
          3378 => x"7e", -- $00d32
          3379 => x"7d", -- $00d33
          3380 => x"7d", -- $00d34
          3381 => x"7d", -- $00d35
          3382 => x"7d", -- $00d36
          3383 => x"7d", -- $00d37
          3384 => x"7d", -- $00d38
          3385 => x"7c", -- $00d39
          3386 => x"7d", -- $00d3a
          3387 => x"7e", -- $00d3b
          3388 => x"7c", -- $00d3c
          3389 => x"7d", -- $00d3d
          3390 => x"7d", -- $00d3e
          3391 => x"7d", -- $00d3f
          3392 => x"7d", -- $00d40
          3393 => x"7d", -- $00d41
          3394 => x"7d", -- $00d42
          3395 => x"7c", -- $00d43
          3396 => x"7d", -- $00d44
          3397 => x"7d", -- $00d45
          3398 => x"7d", -- $00d46
          3399 => x"7c", -- $00d47
          3400 => x"7d", -- $00d48
          3401 => x"7e", -- $00d49
          3402 => x"7d", -- $00d4a
          3403 => x"7d", -- $00d4b
          3404 => x"7d", -- $00d4c
          3405 => x"7d", -- $00d4d
          3406 => x"7d", -- $00d4e
          3407 => x"7d", -- $00d4f
          3408 => x"7d", -- $00d50
          3409 => x"7d", -- $00d51
          3410 => x"7e", -- $00d52
          3411 => x"7d", -- $00d53
          3412 => x"7d", -- $00d54
          3413 => x"7d", -- $00d55
          3414 => x"7d", -- $00d56
          3415 => x"7d", -- $00d57
          3416 => x"7d", -- $00d58
          3417 => x"7d", -- $00d59
          3418 => x"7d", -- $00d5a
          3419 => x"7d", -- $00d5b
          3420 => x"7d", -- $00d5c
          3421 => x"7d", -- $00d5d
          3422 => x"7d", -- $00d5e
          3423 => x"7d", -- $00d5f
          3424 => x"7d", -- $00d60
          3425 => x"7d", -- $00d61
          3426 => x"7d", -- $00d62
          3427 => x"7d", -- $00d63
          3428 => x"7d", -- $00d64
          3429 => x"7e", -- $00d65
          3430 => x"7d", -- $00d66
          3431 => x"7d", -- $00d67
          3432 => x"7d", -- $00d68
          3433 => x"7e", -- $00d69
          3434 => x"7d", -- $00d6a
          3435 => x"7d", -- $00d6b
          3436 => x"7d", -- $00d6c
          3437 => x"7d", -- $00d6d
          3438 => x"7e", -- $00d6e
          3439 => x"7d", -- $00d6f
          3440 => x"7d", -- $00d70
          3441 => x"7d", -- $00d71
          3442 => x"7e", -- $00d72
          3443 => x"7e", -- $00d73
          3444 => x"7e", -- $00d74
          3445 => x"7d", -- $00d75
          3446 => x"7e", -- $00d76
          3447 => x"7e", -- $00d77
          3448 => x"7e", -- $00d78
          3449 => x"7e", -- $00d79
          3450 => x"7d", -- $00d7a
          3451 => x"7e", -- $00d7b
          3452 => x"7e", -- $00d7c
          3453 => x"7e", -- $00d7d
          3454 => x"7d", -- $00d7e
          3455 => x"7e", -- $00d7f
          3456 => x"7e", -- $00d80
          3457 => x"7e", -- $00d81
          3458 => x"7d", -- $00d82
          3459 => x"7d", -- $00d83
          3460 => x"7e", -- $00d84
          3461 => x"7e", -- $00d85
          3462 => x"7e", -- $00d86
          3463 => x"7d", -- $00d87
          3464 => x"7e", -- $00d88
          3465 => x"7e", -- $00d89
          3466 => x"7e", -- $00d8a
          3467 => x"7e", -- $00d8b
          3468 => x"7e", -- $00d8c
          3469 => x"7e", -- $00d8d
          3470 => x"7e", -- $00d8e
          3471 => x"7e", -- $00d8f
          3472 => x"7e", -- $00d90
          3473 => x"7e", -- $00d91
          3474 => x"7e", -- $00d92
          3475 => x"7e", -- $00d93
          3476 => x"7d", -- $00d94
          3477 => x"7d", -- $00d95
          3478 => x"7e", -- $00d96
          3479 => x"7e", -- $00d97
          3480 => x"7e", -- $00d98
          3481 => x"7d", -- $00d99
          3482 => x"7e", -- $00d9a
          3483 => x"7e", -- $00d9b
          3484 => x"7e", -- $00d9c
          3485 => x"7e", -- $00d9d
          3486 => x"7e", -- $00d9e
          3487 => x"7e", -- $00d9f
          3488 => x"7e", -- $00da0
          3489 => x"7e", -- $00da1
          3490 => x"7e", -- $00da2
          3491 => x"7e", -- $00da3
          3492 => x"7e", -- $00da4
          3493 => x"7e", -- $00da5
          3494 => x"7e", -- $00da6
          3495 => x"7e", -- $00da7
          3496 => x"7e", -- $00da8
          3497 => x"7e", -- $00da9
          3498 => x"7e", -- $00daa
          3499 => x"7e", -- $00dab
          3500 => x"7e", -- $00dac
          3501 => x"7e", -- $00dad
          3502 => x"7e", -- $00dae
          3503 => x"7e", -- $00daf
          3504 => x"7e", -- $00db0
          3505 => x"7e", -- $00db1
          3506 => x"7e", -- $00db2
          3507 => x"7e", -- $00db3
          3508 => x"7e", -- $00db4
          3509 => x"7e", -- $00db5
          3510 => x"7e", -- $00db6
          3511 => x"7e", -- $00db7
          3512 => x"7e", -- $00db8
          3513 => x"7e", -- $00db9
          3514 => x"7e", -- $00dba
          3515 => x"7e", -- $00dbb
          3516 => x"7e", -- $00dbc
          3517 => x"7e", -- $00dbd
          3518 => x"7e", -- $00dbe
          3519 => x"7e", -- $00dbf
          3520 => x"7e", -- $00dc0
          3521 => x"7e", -- $00dc1
          3522 => x"7f", -- $00dc2
          3523 => x"7f", -- $00dc3
          3524 => x"7f", -- $00dc4
          3525 => x"7f", -- $00dc5
          3526 => x"7f", -- $00dc6
          3527 => x"7f", -- $00dc7
          3528 => x"7f", -- $00dc8
          3529 => x"7f", -- $00dc9
          3530 => x"7f", -- $00dca
          3531 => x"7f", -- $00dcb
          3532 => x"7f", -- $00dcc
          3533 => x"7f", -- $00dcd
          3534 => x"7f", -- $00dce
          3535 => x"7f", -- $00dcf
          3536 => x"7f", -- $00dd0
          3537 => x"7f", -- $00dd1
          3538 => x"7f", -- $00dd2
          3539 => x"7f", -- $00dd3
          3540 => x"7f", -- $00dd4
          3541 => x"7f", -- $00dd5
          3542 => x"7f", -- $00dd6
          3543 => x"7f", -- $00dd7
          3544 => x"7f", -- $00dd8
          3545 => x"7f", -- $00dd9
          3546 => x"7f", -- $00dda
          3547 => x"7f", -- $00ddb
          3548 => x"7f", -- $00ddc
          3549 => x"7f", -- $00ddd
          3550 => x"7f", -- $00dde
          3551 => x"7f", -- $00ddf
          3552 => x"7f", -- $00de0
          3553 => x"7f", -- $00de1
          3554 => x"7f", -- $00de2
          3555 => x"7f", -- $00de3
          3556 => x"7f", -- $00de4
          3557 => x"80", -- $00de5
          3558 => x"7f", -- $00de6
          3559 => x"80", -- $00de7
          3560 => x"80", -- $00de8
          3561 => x"80", -- $00de9
          3562 => x"80", -- $00dea
          3563 => x"80", -- $00deb
          3564 => x"80", -- $00dec
          3565 => x"80", -- $00ded
          3566 => x"80", -- $00dee
          3567 => x"80", -- $00def
          3568 => x"80", -- $00df0
          3569 => x"80", -- $00df1
          3570 => x"80", -- $00df2
          3571 => x"80", -- $00df3
          3572 => x"80", -- $00df4
          3573 => x"80", -- $00df5
          3574 => x"80", -- $00df6
          3575 => x"80", -- $00df7
          3576 => x"80", -- $00df8
          3577 => x"80", -- $00df9
          3578 => x"80", -- $00dfa
          3579 => x"80", -- $00dfb
          3580 => x"80", -- $00dfc
          3581 => x"80", -- $00dfd
          3582 => x"80", -- $00dfe
          3583 => x"80", -- $00dff
          3584 => x"80", -- $00e00
          3585 => x"80", -- $00e01
          3586 => x"80", -- $00e02
          3587 => x"80", -- $00e03
          3588 => x"80", -- $00e04
          3589 => x"80", -- $00e05
          3590 => x"80", -- $00e06
          3591 => x"80", -- $00e07
          3592 => x"80", -- $00e08
          3593 => x"80", -- $00e09
          3594 => x"80", -- $00e0a
          3595 => x"80", -- $00e0b
          3596 => x"80", -- $00e0c
          3597 => x"80", -- $00e0d
          3598 => x"80", -- $00e0e
          3599 => x"80", -- $00e0f
          3600 => x"80", -- $00e10
          3601 => x"80", -- $00e11
          3602 => x"80", -- $00e12
          3603 => x"80", -- $00e13
          3604 => x"80", -- $00e14
          3605 => x"80", -- $00e15
          3606 => x"80", -- $00e16
          3607 => x"80", -- $00e17
          3608 => x"80", -- $00e18
          3609 => x"80", -- $00e19
          3610 => x"80", -- $00e1a
          3611 => x"80", -- $00e1b
          3612 => x"80", -- $00e1c
          3613 => x"80", -- $00e1d
          3614 => x"81", -- $00e1e
          3615 => x"81", -- $00e1f
          3616 => x"81", -- $00e20
          3617 => x"81", -- $00e21
          3618 => x"81", -- $00e22
          3619 => x"81", -- $00e23
          3620 => x"81", -- $00e24
          3621 => x"81", -- $00e25
          3622 => x"81", -- $00e26
          3623 => x"81", -- $00e27
          3624 => x"81", -- $00e28
          3625 => x"81", -- $00e29
          3626 => x"81", -- $00e2a
          3627 => x"81", -- $00e2b
          3628 => x"81", -- $00e2c
          3629 => x"81", -- $00e2d
          3630 => x"81", -- $00e2e
          3631 => x"81", -- $00e2f
          3632 => x"81", -- $00e30
          3633 => x"81", -- $00e31
          3634 => x"81", -- $00e32
          3635 => x"81", -- $00e33
          3636 => x"81", -- $00e34
          3637 => x"82", -- $00e35
          3638 => x"82", -- $00e36
          3639 => x"82", -- $00e37
          3640 => x"81", -- $00e38
          3641 => x"82", -- $00e39
          3642 => x"82", -- $00e3a
          3643 => x"82", -- $00e3b
          3644 => x"81", -- $00e3c
          3645 => x"82", -- $00e3d
          3646 => x"82", -- $00e3e
          3647 => x"82", -- $00e3f
          3648 => x"82", -- $00e40
          3649 => x"82", -- $00e41
          3650 => x"82", -- $00e42
          3651 => x"82", -- $00e43
          3652 => x"82", -- $00e44
          3653 => x"82", -- $00e45
          3654 => x"82", -- $00e46
          3655 => x"82", -- $00e47
          3656 => x"83", -- $00e48
          3657 => x"82", -- $00e49
          3658 => x"82", -- $00e4a
          3659 => x"82", -- $00e4b
          3660 => x"82", -- $00e4c
          3661 => x"82", -- $00e4d
          3662 => x"82", -- $00e4e
          3663 => x"83", -- $00e4f
          3664 => x"83", -- $00e50
          3665 => x"83", -- $00e51
          3666 => x"83", -- $00e52
          3667 => x"83", -- $00e53
          3668 => x"83", -- $00e54
          3669 => x"82", -- $00e55
          3670 => x"83", -- $00e56
          3671 => x"83", -- $00e57
          3672 => x"83", -- $00e58
          3673 => x"82", -- $00e59
          3674 => x"82", -- $00e5a
          3675 => x"83", -- $00e5b
          3676 => x"83", -- $00e5c
          3677 => x"83", -- $00e5d
          3678 => x"83", -- $00e5e
          3679 => x"83", -- $00e5f
          3680 => x"83", -- $00e60
          3681 => x"83", -- $00e61
          3682 => x"83", -- $00e62
          3683 => x"83", -- $00e63
          3684 => x"83", -- $00e64
          3685 => x"83", -- $00e65
          3686 => x"83", -- $00e66
          3687 => x"83", -- $00e67
          3688 => x"83", -- $00e68
          3689 => x"83", -- $00e69
          3690 => x"83", -- $00e6a
          3691 => x"83", -- $00e6b
          3692 => x"83", -- $00e6c
          3693 => x"83", -- $00e6d
          3694 => x"83", -- $00e6e
          3695 => x"83", -- $00e6f
          3696 => x"83", -- $00e70
          3697 => x"83", -- $00e71
          3698 => x"83", -- $00e72
          3699 => x"83", -- $00e73
          3700 => x"83", -- $00e74
          3701 => x"83", -- $00e75
          3702 => x"83", -- $00e76
          3703 => x"83", -- $00e77
          3704 => x"83", -- $00e78
          3705 => x"83", -- $00e79
          3706 => x"83", -- $00e7a
          3707 => x"83", -- $00e7b
          3708 => x"83", -- $00e7c
          3709 => x"82", -- $00e7d
          3710 => x"82", -- $00e7e
          3711 => x"83", -- $00e7f
          3712 => x"83", -- $00e80
          3713 => x"82", -- $00e81
          3714 => x"82", -- $00e82
          3715 => x"83", -- $00e83
          3716 => x"83", -- $00e84
          3717 => x"83", -- $00e85
          3718 => x"83", -- $00e86
          3719 => x"83", -- $00e87
          3720 => x"83", -- $00e88
          3721 => x"83", -- $00e89
          3722 => x"82", -- $00e8a
          3723 => x"82", -- $00e8b
          3724 => x"83", -- $00e8c
          3725 => x"83", -- $00e8d
          3726 => x"82", -- $00e8e
          3727 => x"82", -- $00e8f
          3728 => x"82", -- $00e90
          3729 => x"82", -- $00e91
          3730 => x"82", -- $00e92
          3731 => x"82", -- $00e93
          3732 => x"82", -- $00e94
          3733 => x"82", -- $00e95
          3734 => x"82", -- $00e96
          3735 => x"82", -- $00e97
          3736 => x"82", -- $00e98
          3737 => x"82", -- $00e99
          3738 => x"82", -- $00e9a
          3739 => x"82", -- $00e9b
          3740 => x"82", -- $00e9c
          3741 => x"82", -- $00e9d
          3742 => x"82", -- $00e9e
          3743 => x"82", -- $00e9f
          3744 => x"82", -- $00ea0
          3745 => x"82", -- $00ea1
          3746 => x"82", -- $00ea2
          3747 => x"82", -- $00ea3
          3748 => x"82", -- $00ea4
          3749 => x"82", -- $00ea5
          3750 => x"82", -- $00ea6
          3751 => x"83", -- $00ea7
          3752 => x"83", -- $00ea8
          3753 => x"83", -- $00ea9
          3754 => x"83", -- $00eaa
          3755 => x"83", -- $00eab
          3756 => x"83", -- $00eac
          3757 => x"82", -- $00ead
          3758 => x"83", -- $00eae
          3759 => x"83", -- $00eaf
          3760 => x"83", -- $00eb0
          3761 => x"82", -- $00eb1
          3762 => x"83", -- $00eb2
          3763 => x"83", -- $00eb3
          3764 => x"83", -- $00eb4
          3765 => x"82", -- $00eb5
          3766 => x"82", -- $00eb6
          3767 => x"83", -- $00eb7
          3768 => x"83", -- $00eb8
          3769 => x"83", -- $00eb9
          3770 => x"83", -- $00eba
          3771 => x"83", -- $00ebb
          3772 => x"83", -- $00ebc
          3773 => x"83", -- $00ebd
          3774 => x"83", -- $00ebe
          3775 => x"83", -- $00ebf
          3776 => x"83", -- $00ec0
          3777 => x"83", -- $00ec1
          3778 => x"83", -- $00ec2
          3779 => x"83", -- $00ec3
          3780 => x"83", -- $00ec4
          3781 => x"83", -- $00ec5
          3782 => x"83", -- $00ec6
          3783 => x"83", -- $00ec7
          3784 => x"83", -- $00ec8
          3785 => x"83", -- $00ec9
          3786 => x"84", -- $00eca
          3787 => x"84", -- $00ecb
          3788 => x"83", -- $00ecc
          3789 => x"83", -- $00ecd
          3790 => x"83", -- $00ece
          3791 => x"84", -- $00ecf
          3792 => x"83", -- $00ed0
          3793 => x"83", -- $00ed1
          3794 => x"83", -- $00ed2
          3795 => x"83", -- $00ed3
          3796 => x"84", -- $00ed4
          3797 => x"83", -- $00ed5
          3798 => x"83", -- $00ed6
          3799 => x"83", -- $00ed7
          3800 => x"83", -- $00ed8
          3801 => x"83", -- $00ed9
          3802 => x"83", -- $00eda
          3803 => x"83", -- $00edb
          3804 => x"83", -- $00edc
          3805 => x"83", -- $00edd
          3806 => x"83", -- $00ede
          3807 => x"83", -- $00edf
          3808 => x"83", -- $00ee0
          3809 => x"84", -- $00ee1
          3810 => x"84", -- $00ee2
          3811 => x"83", -- $00ee3
          3812 => x"83", -- $00ee4
          3813 => x"83", -- $00ee5
          3814 => x"83", -- $00ee6
          3815 => x"83", -- $00ee7
          3816 => x"83", -- $00ee8
          3817 => x"83", -- $00ee9
          3818 => x"83", -- $00eea
          3819 => x"83", -- $00eeb
          3820 => x"83", -- $00eec
          3821 => x"83", -- $00eed
          3822 => x"83", -- $00eee
          3823 => x"83", -- $00eef
          3824 => x"83", -- $00ef0
          3825 => x"83", -- $00ef1
          3826 => x"83", -- $00ef2
          3827 => x"83", -- $00ef3
          3828 => x"83", -- $00ef4
          3829 => x"83", -- $00ef5
          3830 => x"83", -- $00ef6
          3831 => x"83", -- $00ef7
          3832 => x"83", -- $00ef8
          3833 => x"83", -- $00ef9
          3834 => x"83", -- $00efa
          3835 => x"83", -- $00efb
          3836 => x"83", -- $00efc
          3837 => x"83", -- $00efd
          3838 => x"83", -- $00efe
          3839 => x"83", -- $00eff
          3840 => x"83", -- $00f00
          3841 => x"83", -- $00f01
          3842 => x"83", -- $00f02
          3843 => x"83", -- $00f03
          3844 => x"83", -- $00f04
          3845 => x"83", -- $00f05
          3846 => x"83", -- $00f06
          3847 => x"83", -- $00f07
          3848 => x"83", -- $00f08
          3849 => x"83", -- $00f09
          3850 => x"83", -- $00f0a
          3851 => x"83", -- $00f0b
          3852 => x"82", -- $00f0c
          3853 => x"82", -- $00f0d
          3854 => x"82", -- $00f0e
          3855 => x"82", -- $00f0f
          3856 => x"82", -- $00f10
          3857 => x"82", -- $00f11
          3858 => x"82", -- $00f12
          3859 => x"82", -- $00f13
          3860 => x"82", -- $00f14
          3861 => x"82", -- $00f15
          3862 => x"82", -- $00f16
          3863 => x"82", -- $00f17
          3864 => x"82", -- $00f18
          3865 => x"82", -- $00f19
          3866 => x"82", -- $00f1a
          3867 => x"82", -- $00f1b
          3868 => x"82", -- $00f1c
          3869 => x"82", -- $00f1d
          3870 => x"82", -- $00f1e
          3871 => x"82", -- $00f1f
          3872 => x"82", -- $00f20
          3873 => x"82", -- $00f21
          3874 => x"82", -- $00f22
          3875 => x"82", -- $00f23
          3876 => x"82", -- $00f24
          3877 => x"82", -- $00f25
          3878 => x"82", -- $00f26
          3879 => x"82", -- $00f27
          3880 => x"82", -- $00f28
          3881 => x"82", -- $00f29
          3882 => x"82", -- $00f2a
          3883 => x"82", -- $00f2b
          3884 => x"82", -- $00f2c
          3885 => x"82", -- $00f2d
          3886 => x"82", -- $00f2e
          3887 => x"82", -- $00f2f
          3888 => x"82", -- $00f30
          3889 => x"82", -- $00f31
          3890 => x"82", -- $00f32
          3891 => x"82", -- $00f33
          3892 => x"82", -- $00f34
          3893 => x"82", -- $00f35
          3894 => x"82", -- $00f36
          3895 => x"82", -- $00f37
          3896 => x"81", -- $00f38
          3897 => x"82", -- $00f39
          3898 => x"82", -- $00f3a
          3899 => x"81", -- $00f3b
          3900 => x"81", -- $00f3c
          3901 => x"81", -- $00f3d
          3902 => x"81", -- $00f3e
          3903 => x"81", -- $00f3f
          3904 => x"81", -- $00f40
          3905 => x"81", -- $00f41
          3906 => x"81", -- $00f42
          3907 => x"81", -- $00f43
          3908 => x"81", -- $00f44
          3909 => x"81", -- $00f45
          3910 => x"81", -- $00f46
          3911 => x"81", -- $00f47
          3912 => x"81", -- $00f48
          3913 => x"81", -- $00f49
          3914 => x"81", -- $00f4a
          3915 => x"81", -- $00f4b
          3916 => x"81", -- $00f4c
          3917 => x"81", -- $00f4d
          3918 => x"81", -- $00f4e
          3919 => x"81", -- $00f4f
          3920 => x"81", -- $00f50
          3921 => x"81", -- $00f51
          3922 => x"81", -- $00f52
          3923 => x"81", -- $00f53
          3924 => x"81", -- $00f54
          3925 => x"81", -- $00f55
          3926 => x"81", -- $00f56
          3927 => x"81", -- $00f57
          3928 => x"81", -- $00f58
          3929 => x"81", -- $00f59
          3930 => x"81", -- $00f5a
          3931 => x"81", -- $00f5b
          3932 => x"81", -- $00f5c
          3933 => x"81", -- $00f5d
          3934 => x"80", -- $00f5e
          3935 => x"80", -- $00f5f
          3936 => x"80", -- $00f60
          3937 => x"80", -- $00f61
          3938 => x"80", -- $00f62
          3939 => x"80", -- $00f63
          3940 => x"80", -- $00f64
          3941 => x"80", -- $00f65
          3942 => x"80", -- $00f66
          3943 => x"80", -- $00f67
          3944 => x"80", -- $00f68
          3945 => x"80", -- $00f69
          3946 => x"80", -- $00f6a
          3947 => x"80", -- $00f6b
          3948 => x"80", -- $00f6c
          3949 => x"80", -- $00f6d
          3950 => x"80", -- $00f6e
          3951 => x"80", -- $00f6f
          3952 => x"80", -- $00f70
          3953 => x"80", -- $00f71
          3954 => x"80", -- $00f72
          3955 => x"80", -- $00f73
          3956 => x"80", -- $00f74
          3957 => x"80", -- $00f75
          3958 => x"80", -- $00f76
          3959 => x"80", -- $00f77
          3960 => x"80", -- $00f78
          3961 => x"80", -- $00f79
          3962 => x"80", -- $00f7a
          3963 => x"80", -- $00f7b
          3964 => x"80", -- $00f7c
          3965 => x"80", -- $00f7d
          3966 => x"80", -- $00f7e
          3967 => x"80", -- $00f7f
          3968 => x"80", -- $00f80
          3969 => x"80", -- $00f81
          3970 => x"80", -- $00f82
          3971 => x"80", -- $00f83
          3972 => x"80", -- $00f84
          3973 => x"80", -- $00f85
          3974 => x"80", -- $00f86
          3975 => x"80", -- $00f87
          3976 => x"7f", -- $00f88
          3977 => x"7f", -- $00f89
          3978 => x"7f", -- $00f8a
          3979 => x"7f", -- $00f8b
          3980 => x"7f", -- $00f8c
          3981 => x"7f", -- $00f8d
          3982 => x"7f", -- $00f8e
          3983 => x"7f", -- $00f8f
          3984 => x"7f", -- $00f90
          3985 => x"7f", -- $00f91
          3986 => x"7f", -- $00f92
          3987 => x"7f", -- $00f93
          3988 => x"7f", -- $00f94
          3989 => x"7f", -- $00f95
          3990 => x"7f", -- $00f96
          3991 => x"7f", -- $00f97
          3992 => x"7f", -- $00f98
          3993 => x"7f", -- $00f99
          3994 => x"7f", -- $00f9a
          3995 => x"7f", -- $00f9b
          3996 => x"7f", -- $00f9c
          3997 => x"7f", -- $00f9d
          3998 => x"7f", -- $00f9e
          3999 => x"7f", -- $00f9f
          4000 => x"7f", -- $00fa0
          4001 => x"7f", -- $00fa1
          4002 => x"7f", -- $00fa2
          4003 => x"7f", -- $00fa3
          4004 => x"7f", -- $00fa4
          4005 => x"7f", -- $00fa5
          4006 => x"7f", -- $00fa6
          4007 => x"7f", -- $00fa7
          4008 => x"7f", -- $00fa8
          4009 => x"7f", -- $00fa9
          4010 => x"7f", -- $00faa
          4011 => x"7e", -- $00fab
          4012 => x"7e", -- $00fac
          4013 => x"7e", -- $00fad
          4014 => x"7e", -- $00fae
          4015 => x"7e", -- $00faf
          4016 => x"7e", -- $00fb0
          4017 => x"7e", -- $00fb1
          4018 => x"7e", -- $00fb2
          4019 => x"7e", -- $00fb3
          4020 => x"7e", -- $00fb4
          4021 => x"7e", -- $00fb5
          4022 => x"7e", -- $00fb6
          4023 => x"7e", -- $00fb7
          4024 => x"7e", -- $00fb8
          4025 => x"7e", -- $00fb9
          4026 => x"7e", -- $00fba
          4027 => x"7e", -- $00fbb
          4028 => x"7e", -- $00fbc
          4029 => x"7e", -- $00fbd
          4030 => x"7e", -- $00fbe
          4031 => x"7e", -- $00fbf
          4032 => x"7e", -- $00fc0
          4033 => x"7e", -- $00fc1
          4034 => x"7e", -- $00fc2
          4035 => x"7e", -- $00fc3
          4036 => x"7e", -- $00fc4
          4037 => x"7e", -- $00fc5
          4038 => x"7e", -- $00fc6
          4039 => x"7e", -- $00fc7
          4040 => x"7e", -- $00fc8
          4041 => x"7e", -- $00fc9
          4042 => x"7e", -- $00fca
          4043 => x"7e", -- $00fcb
          4044 => x"7e", -- $00fcc
          4045 => x"7d", -- $00fcd
          4046 => x"7e", -- $00fce
          4047 => x"7e", -- $00fcf
          4048 => x"7e", -- $00fd0
          4049 => x"7e", -- $00fd1
          4050 => x"7d", -- $00fd2
          4051 => x"7d", -- $00fd3
          4052 => x"7d", -- $00fd4
          4053 => x"7d", -- $00fd5
          4054 => x"7d", -- $00fd6
          4055 => x"7d", -- $00fd7
          4056 => x"7d", -- $00fd8
          4057 => x"7d", -- $00fd9
          4058 => x"7d", -- $00fda
          4059 => x"7d", -- $00fdb
          4060 => x"7d", -- $00fdc
          4061 => x"7d", -- $00fdd
          4062 => x"7d", -- $00fde
          4063 => x"7d", -- $00fdf
          4064 => x"7d", -- $00fe0
          4065 => x"7d", -- $00fe1
          4066 => x"7d", -- $00fe2
          4067 => x"7d", -- $00fe3
          4068 => x"7d", -- $00fe4
          4069 => x"7d", -- $00fe5
          4070 => x"7d", -- $00fe6
          4071 => x"7d", -- $00fe7
          4072 => x"7e", -- $00fe8
          4073 => x"7e", -- $00fe9
          4074 => x"7d", -- $00fea
          4075 => x"7d", -- $00feb
          4076 => x"7d", -- $00fec
          4077 => x"7d", -- $00fed
          4078 => x"7d", -- $00fee
          4079 => x"7d", -- $00fef
          4080 => x"7d", -- $00ff0
          4081 => x"7d", -- $00ff1
          4082 => x"7d", -- $00ff2
          4083 => x"7d", -- $00ff3
          4084 => x"7d", -- $00ff4
          4085 => x"7d", -- $00ff5
          4086 => x"7d", -- $00ff6
          4087 => x"7d", -- $00ff7
          4088 => x"7d", -- $00ff8
          4089 => x"7d", -- $00ff9
          4090 => x"7d", -- $00ffa
          4091 => x"7d", -- $00ffb
          4092 => x"7d", -- $00ffc
          4093 => x"7d", -- $00ffd
          4094 => x"7d", -- $00ffe
          4095 => x"7d", -- $00fff
          4096 => x"7d", -- $01000
          4097 => x"7d", -- $01001
          4098 => x"7d", -- $01002
          4099 => x"7d", -- $01003
          4100 => x"7d", -- $01004
          4101 => x"7d", -- $01005
          4102 => x"7d", -- $01006
          4103 => x"7d", -- $01007
          4104 => x"7d", -- $01008
          4105 => x"7d", -- $01009
          4106 => x"7d", -- $0100a
          4107 => x"7d", -- $0100b
          4108 => x"7d", -- $0100c
          4109 => x"7d", -- $0100d
          4110 => x"7d", -- $0100e
          4111 => x"7d", -- $0100f
          4112 => x"7d", -- $01010
          4113 => x"7d", -- $01011
          4114 => x"7d", -- $01012
          4115 => x"7d", -- $01013
          4116 => x"7d", -- $01014
          4117 => x"7d", -- $01015
          4118 => x"7d", -- $01016
          4119 => x"7d", -- $01017
          4120 => x"7d", -- $01018
          4121 => x"7d", -- $01019
          4122 => x"7d", -- $0101a
          4123 => x"7d", -- $0101b
          4124 => x"7d", -- $0101c
          4125 => x"7d", -- $0101d
          4126 => x"7d", -- $0101e
          4127 => x"7d", -- $0101f
          4128 => x"7d", -- $01020
          4129 => x"7d", -- $01021
          4130 => x"7d", -- $01022
          4131 => x"7d", -- $01023
          4132 => x"7d", -- $01024
          4133 => x"7d", -- $01025
          4134 => x"7d", -- $01026
          4135 => x"7d", -- $01027
          4136 => x"7d", -- $01028
          4137 => x"7d", -- $01029
          4138 => x"7d", -- $0102a
          4139 => x"7d", -- $0102b
          4140 => x"7d", -- $0102c
          4141 => x"7d", -- $0102d
          4142 => x"7c", -- $0102e
          4143 => x"7c", -- $0102f
          4144 => x"7c", -- $01030
          4145 => x"7c", -- $01031
          4146 => x"7d", -- $01032
          4147 => x"7d", -- $01033
          4148 => x"7c", -- $01034
          4149 => x"7d", -- $01035
          4150 => x"7c", -- $01036
          4151 => x"7c", -- $01037
          4152 => x"7c", -- $01038
          4153 => x"7c", -- $01039
          4154 => x"7c", -- $0103a
          4155 => x"7c", -- $0103b
          4156 => x"7c", -- $0103c
          4157 => x"7c", -- $0103d
          4158 => x"7c", -- $0103e
          4159 => x"7c", -- $0103f
          4160 => x"7c", -- $01040
          4161 => x"7c", -- $01041
          4162 => x"7c", -- $01042
          4163 => x"7c", -- $01043
          4164 => x"7c", -- $01044
          4165 => x"7c", -- $01045
          4166 => x"7c", -- $01046
          4167 => x"7c", -- $01047
          4168 => x"7c", -- $01048
          4169 => x"7c", -- $01049
          4170 => x"7c", -- $0104a
          4171 => x"7c", -- $0104b
          4172 => x"7c", -- $0104c
          4173 => x"7c", -- $0104d
          4174 => x"7c", -- $0104e
          4175 => x"7c", -- $0104f
          4176 => x"7c", -- $01050
          4177 => x"7c", -- $01051
          4178 => x"7c", -- $01052
          4179 => x"7c", -- $01053
          4180 => x"7c", -- $01054
          4181 => x"7c", -- $01055
          4182 => x"7c", -- $01056
          4183 => x"7c", -- $01057
          4184 => x"7c", -- $01058
          4185 => x"7c", -- $01059
          4186 => x"7c", -- $0105a
          4187 => x"7c", -- $0105b
          4188 => x"7c", -- $0105c
          4189 => x"7c", -- $0105d
          4190 => x"7c", -- $0105e
          4191 => x"7c", -- $0105f
          4192 => x"7c", -- $01060
          4193 => x"7c", -- $01061
          4194 => x"7c", -- $01062
          4195 => x"7c", -- $01063
          4196 => x"7c", -- $01064
          4197 => x"7c", -- $01065
          4198 => x"7c", -- $01066
          4199 => x"7c", -- $01067
          4200 => x"7c", -- $01068
          4201 => x"7c", -- $01069
          4202 => x"7d", -- $0106a
          4203 => x"7d", -- $0106b
          4204 => x"7d", -- $0106c
          4205 => x"7d", -- $0106d
          4206 => x"7d", -- $0106e
          4207 => x"7d", -- $0106f
          4208 => x"7d", -- $01070
          4209 => x"7d", -- $01071
          4210 => x"7d", -- $01072
          4211 => x"7d", -- $01073
          4212 => x"7d", -- $01074
          4213 => x"7d", -- $01075
          4214 => x"7d", -- $01076
          4215 => x"7d", -- $01077
          4216 => x"7d", -- $01078
          4217 => x"7d", -- $01079
          4218 => x"7d", -- $0107a
          4219 => x"7d", -- $0107b
          4220 => x"7d", -- $0107c
          4221 => x"7d", -- $0107d
          4222 => x"7d", -- $0107e
          4223 => x"7d", -- $0107f
          4224 => x"7d", -- $01080
          4225 => x"7d", -- $01081
          4226 => x"7d", -- $01082
          4227 => x"7d", -- $01083
          4228 => x"7d", -- $01084
          4229 => x"7d", -- $01085
          4230 => x"7d", -- $01086
          4231 => x"7d", -- $01087
          4232 => x"7d", -- $01088
          4233 => x"7d", -- $01089
          4234 => x"7d", -- $0108a
          4235 => x"7d", -- $0108b
          4236 => x"7d", -- $0108c
          4237 => x"7d", -- $0108d
          4238 => x"7d", -- $0108e
          4239 => x"7d", -- $0108f
          4240 => x"7e", -- $01090
          4241 => x"7e", -- $01091
          4242 => x"7e", -- $01092
          4243 => x"7e", -- $01093
          4244 => x"7e", -- $01094
          4245 => x"7e", -- $01095
          4246 => x"7e", -- $01096
          4247 => x"7e", -- $01097
          4248 => x"7e", -- $01098
          4249 => x"7e", -- $01099
          4250 => x"7e", -- $0109a
          4251 => x"7e", -- $0109b
          4252 => x"7e", -- $0109c
          4253 => x"7e", -- $0109d
          4254 => x"7e", -- $0109e
          4255 => x"7e", -- $0109f
          4256 => x"7e", -- $010a0
          4257 => x"7e", -- $010a1
          4258 => x"7e", -- $010a2
          4259 => x"7e", -- $010a3
          4260 => x"7e", -- $010a4
          4261 => x"7e", -- $010a5
          4262 => x"7e", -- $010a6
          4263 => x"7e", -- $010a7
          4264 => x"7e", -- $010a8
          4265 => x"7f", -- $010a9
          4266 => x"7f", -- $010aa
          4267 => x"7f", -- $010ab
          4268 => x"7f", -- $010ac
          4269 => x"7f", -- $010ad
          4270 => x"7f", -- $010ae
          4271 => x"7f", -- $010af
          4272 => x"7f", -- $010b0
          4273 => x"7f", -- $010b1
          4274 => x"7f", -- $010b2
          4275 => x"7f", -- $010b3
          4276 => x"7f", -- $010b4
          4277 => x"7f", -- $010b5
          4278 => x"7f", -- $010b6
          4279 => x"7f", -- $010b7
          4280 => x"7f", -- $010b8
          4281 => x"7f", -- $010b9
          4282 => x"7f", -- $010ba
          4283 => x"7f", -- $010bb
          4284 => x"7f", -- $010bc
          4285 => x"7f", -- $010bd
          4286 => x"7f", -- $010be
          4287 => x"7f", -- $010bf
          4288 => x"7f", -- $010c0
          4289 => x"7f", -- $010c1
          4290 => x"80", -- $010c2
          4291 => x"7f", -- $010c3
          4292 => x"7f", -- $010c4
          4293 => x"7f", -- $010c5
          4294 => x"80", -- $010c6
          4295 => x"80", -- $010c7
          4296 => x"80", -- $010c8
          4297 => x"80", -- $010c9
          4298 => x"7f", -- $010ca
          4299 => x"7f", -- $010cb
          4300 => x"7f", -- $010cc
          4301 => x"80", -- $010cd
          4302 => x"80", -- $010ce
          4303 => x"80", -- $010cf
          4304 => x"80", -- $010d0
          4305 => x"80", -- $010d1
          4306 => x"80", -- $010d2
          4307 => x"80", -- $010d3
          4308 => x"80", -- $010d4
          4309 => x"80", -- $010d5
          4310 => x"80", -- $010d6
          4311 => x"80", -- $010d7
          4312 => x"80", -- $010d8
          4313 => x"80", -- $010d9
          4314 => x"80", -- $010da
          4315 => x"80", -- $010db
          4316 => x"80", -- $010dc
          4317 => x"80", -- $010dd
          4318 => x"80", -- $010de
          4319 => x"80", -- $010df
          4320 => x"80", -- $010e0
          4321 => x"80", -- $010e1
          4322 => x"80", -- $010e2
          4323 => x"80", -- $010e3
          4324 => x"80", -- $010e4
          4325 => x"80", -- $010e5
          4326 => x"80", -- $010e6
          4327 => x"80", -- $010e7
          4328 => x"80", -- $010e8
          4329 => x"80", -- $010e9
          4330 => x"80", -- $010ea
          4331 => x"80", -- $010eb
          4332 => x"80", -- $010ec
          4333 => x"80", -- $010ed
          4334 => x"80", -- $010ee
          4335 => x"80", -- $010ef
          4336 => x"80", -- $010f0
          4337 => x"80", -- $010f1
          4338 => x"80", -- $010f2
          4339 => x"80", -- $010f3
          4340 => x"80", -- $010f4
          4341 => x"80", -- $010f5
          4342 => x"80", -- $010f6
          4343 => x"80", -- $010f7
          4344 => x"80", -- $010f8
          4345 => x"80", -- $010f9
          4346 => x"80", -- $010fa
          4347 => x"80", -- $010fb
          4348 => x"80", -- $010fc
          4349 => x"80", -- $010fd
          4350 => x"80", -- $010fe
          4351 => x"80", -- $010ff
          4352 => x"80", -- $01100
          4353 => x"80", -- $01101
          4354 => x"80", -- $01102
          4355 => x"80", -- $01103
          4356 => x"80", -- $01104
          4357 => x"80", -- $01105
          4358 => x"80", -- $01106
          4359 => x"80", -- $01107
          4360 => x"80", -- $01108
          4361 => x"80", -- $01109
          4362 => x"80", -- $0110a
          4363 => x"80", -- $0110b
          4364 => x"80", -- $0110c
          4365 => x"80", -- $0110d
          4366 => x"80", -- $0110e
          4367 => x"80", -- $0110f
          4368 => x"80", -- $01110
          4369 => x"80", -- $01111
          4370 => x"80", -- $01112
          4371 => x"80", -- $01113
          4372 => x"80", -- $01114
          4373 => x"80", -- $01115
          4374 => x"80", -- $01116
          4375 => x"80", -- $01117
          4376 => x"80", -- $01118
          4377 => x"80", -- $01119
          4378 => x"80", -- $0111a
          4379 => x"80", -- $0111b
          4380 => x"80", -- $0111c
          4381 => x"80", -- $0111d
          4382 => x"80", -- $0111e
          4383 => x"80", -- $0111f
          4384 => x"80", -- $01120
          4385 => x"80", -- $01121
          4386 => x"80", -- $01122
          4387 => x"80", -- $01123
          4388 => x"80", -- $01124
          4389 => x"80", -- $01125
          4390 => x"80", -- $01126
          4391 => x"80", -- $01127
          4392 => x"80", -- $01128
          4393 => x"80", -- $01129
          4394 => x"80", -- $0112a
          4395 => x"80", -- $0112b
          4396 => x"80", -- $0112c
          4397 => x"80", -- $0112d
          4398 => x"80", -- $0112e
          4399 => x"80", -- $0112f
          4400 => x"81", -- $01130
          4401 => x"81", -- $01131
          4402 => x"81", -- $01132
          4403 => x"81", -- $01133
          4404 => x"81", -- $01134
          4405 => x"81", -- $01135
          4406 => x"81", -- $01136
          4407 => x"81", -- $01137
          4408 => x"81", -- $01138
          4409 => x"81", -- $01139
          4410 => x"81", -- $0113a
          4411 => x"81", -- $0113b
          4412 => x"81", -- $0113c
          4413 => x"81", -- $0113d
          4414 => x"81", -- $0113e
          4415 => x"81", -- $0113f
          4416 => x"81", -- $01140
          4417 => x"81", -- $01141
          4418 => x"81", -- $01142
          4419 => x"81", -- $01143
          4420 => x"81", -- $01144
          4421 => x"81", -- $01145
          4422 => x"81", -- $01146
          4423 => x"81", -- $01147
          4424 => x"82", -- $01148
          4425 => x"82", -- $01149
          4426 => x"82", -- $0114a
          4427 => x"82", -- $0114b
          4428 => x"81", -- $0114c
          4429 => x"81", -- $0114d
          4430 => x"82", -- $0114e
          4431 => x"81", -- $0114f
          4432 => x"81", -- $01150
          4433 => x"81", -- $01151
          4434 => x"82", -- $01152
          4435 => x"82", -- $01153
          4436 => x"82", -- $01154
          4437 => x"82", -- $01155
          4438 => x"82", -- $01156
          4439 => x"82", -- $01157
          4440 => x"82", -- $01158
          4441 => x"82", -- $01159
          4442 => x"82", -- $0115a
          4443 => x"82", -- $0115b
          4444 => x"82", -- $0115c
          4445 => x"82", -- $0115d
          4446 => x"82", -- $0115e
          4447 => x"82", -- $0115f
          4448 => x"82", -- $01160
          4449 => x"82", -- $01161
          4450 => x"82", -- $01162
          4451 => x"82", -- $01163
          4452 => x"82", -- $01164
          4453 => x"82", -- $01165
          4454 => x"82", -- $01166
          4455 => x"82", -- $01167
          4456 => x"82", -- $01168
          4457 => x"82", -- $01169
          4458 => x"82", -- $0116a
          4459 => x"82", -- $0116b
          4460 => x"82", -- $0116c
          4461 => x"82", -- $0116d
          4462 => x"82", -- $0116e
          4463 => x"82", -- $0116f
          4464 => x"82", -- $01170
          4465 => x"82", -- $01171
          4466 => x"82", -- $01172
          4467 => x"82", -- $01173
          4468 => x"82", -- $01174
          4469 => x"82", -- $01175
          4470 => x"82", -- $01176
          4471 => x"82", -- $01177
          4472 => x"82", -- $01178
          4473 => x"82", -- $01179
          4474 => x"83", -- $0117a
          4475 => x"83", -- $0117b
          4476 => x"83", -- $0117c
          4477 => x"83", -- $0117d
          4478 => x"83", -- $0117e
          4479 => x"83", -- $0117f
          4480 => x"82", -- $01180
          4481 => x"82", -- $01181
          4482 => x"82", -- $01182
          4483 => x"82", -- $01183
          4484 => x"82", -- $01184
          4485 => x"82", -- $01185
          4486 => x"82", -- $01186
          4487 => x"83", -- $01187
          4488 => x"83", -- $01188
          4489 => x"83", -- $01189
          4490 => x"83", -- $0118a
          4491 => x"83", -- $0118b
          4492 => x"83", -- $0118c
          4493 => x"83", -- $0118d
          4494 => x"83", -- $0118e
          4495 => x"83", -- $0118f
          4496 => x"83", -- $01190
          4497 => x"83", -- $01191
          4498 => x"83", -- $01192
          4499 => x"83", -- $01193
          4500 => x"83", -- $01194
          4501 => x"83", -- $01195
          4502 => x"83", -- $01196
          4503 => x"83", -- $01197
          4504 => x"83", -- $01198
          4505 => x"83", -- $01199
          4506 => x"83", -- $0119a
          4507 => x"83", -- $0119b
          4508 => x"83", -- $0119c
          4509 => x"83", -- $0119d
          4510 => x"83", -- $0119e
          4511 => x"83", -- $0119f
          4512 => x"83", -- $011a0
          4513 => x"83", -- $011a1
          4514 => x"83", -- $011a2
          4515 => x"83", -- $011a3
          4516 => x"83", -- $011a4
          4517 => x"83", -- $011a5
          4518 => x"83", -- $011a6
          4519 => x"83", -- $011a7
          4520 => x"83", -- $011a8
          4521 => x"83", -- $011a9
          4522 => x"83", -- $011aa
          4523 => x"83", -- $011ab
          4524 => x"83", -- $011ac
          4525 => x"83", -- $011ad
          4526 => x"83", -- $011ae
          4527 => x"83", -- $011af
          4528 => x"83", -- $011b0
          4529 => x"83", -- $011b1
          4530 => x"83", -- $011b2
          4531 => x"83", -- $011b3
          4532 => x"83", -- $011b4
          4533 => x"83", -- $011b5
          4534 => x"83", -- $011b6
          4535 => x"83", -- $011b7
          4536 => x"83", -- $011b8
          4537 => x"83", -- $011b9
          4538 => x"83", -- $011ba
          4539 => x"83", -- $011bb
          4540 => x"83", -- $011bc
          4541 => x"83", -- $011bd
          4542 => x"83", -- $011be
          4543 => x"83", -- $011bf
          4544 => x"83", -- $011c0
          4545 => x"83", -- $011c1
          4546 => x"83", -- $011c2
          4547 => x"83", -- $011c3
          4548 => x"83", -- $011c4
          4549 => x"83", -- $011c5
          4550 => x"83", -- $011c6
          4551 => x"83", -- $011c7
          4552 => x"83", -- $011c8
          4553 => x"83", -- $011c9
          4554 => x"83", -- $011ca
          4555 => x"83", -- $011cb
          4556 => x"83", -- $011cc
          4557 => x"83", -- $011cd
          4558 => x"83", -- $011ce
          4559 => x"83", -- $011cf
          4560 => x"83", -- $011d0
          4561 => x"83", -- $011d1
          4562 => x"83", -- $011d2
          4563 => x"83", -- $011d3
          4564 => x"83", -- $011d4
          4565 => x"83", -- $011d5
          4566 => x"83", -- $011d6
          4567 => x"83", -- $011d7
          4568 => x"83", -- $011d8
          4569 => x"83", -- $011d9
          4570 => x"83", -- $011da
          4571 => x"83", -- $011db
          4572 => x"83", -- $011dc
          4573 => x"83", -- $011dd
          4574 => x"83", -- $011de
          4575 => x"83", -- $011df
          4576 => x"83", -- $011e0
          4577 => x"83", -- $011e1
          4578 => x"83", -- $011e2
          4579 => x"83", -- $011e3
          4580 => x"83", -- $011e4
          4581 => x"83", -- $011e5
          4582 => x"83", -- $011e6
          4583 => x"83", -- $011e7
          4584 => x"83", -- $011e8
          4585 => x"82", -- $011e9
          4586 => x"82", -- $011ea
          4587 => x"82", -- $011eb
          4588 => x"82", -- $011ec
          4589 => x"82", -- $011ed
          4590 => x"82", -- $011ee
          4591 => x"82", -- $011ef
          4592 => x"82", -- $011f0
          4593 => x"82", -- $011f1
          4594 => x"82", -- $011f2
          4595 => x"82", -- $011f3
          4596 => x"82", -- $011f4
          4597 => x"82", -- $011f5
          4598 => x"82", -- $011f6
          4599 => x"82", -- $011f7
          4600 => x"82", -- $011f8
          4601 => x"82", -- $011f9
          4602 => x"82", -- $011fa
          4603 => x"82", -- $011fb
          4604 => x"82", -- $011fc
          4605 => x"82", -- $011fd
          4606 => x"82", -- $011fe
          4607 => x"82", -- $011ff
          4608 => x"82", -- $01200
          4609 => x"82", -- $01201
          4610 => x"82", -- $01202
          4611 => x"82", -- $01203
          4612 => x"82", -- $01204
          4613 => x"82", -- $01205
          4614 => x"82", -- $01206
          4615 => x"82", -- $01207
          4616 => x"81", -- $01208
          4617 => x"82", -- $01209
          4618 => x"82", -- $0120a
          4619 => x"82", -- $0120b
          4620 => x"82", -- $0120c
          4621 => x"81", -- $0120d
          4622 => x"81", -- $0120e
          4623 => x"81", -- $0120f
          4624 => x"81", -- $01210
          4625 => x"81", -- $01211
          4626 => x"81", -- $01212
          4627 => x"81", -- $01213
          4628 => x"81", -- $01214
          4629 => x"81", -- $01215
          4630 => x"81", -- $01216
          4631 => x"81", -- $01217
          4632 => x"81", -- $01218
          4633 => x"81", -- $01219
          4634 => x"81", -- $0121a
          4635 => x"81", -- $0121b
          4636 => x"81", -- $0121c
          4637 => x"81", -- $0121d
          4638 => x"81", -- $0121e
          4639 => x"81", -- $0121f
          4640 => x"81", -- $01220
          4641 => x"81", -- $01221
          4642 => x"81", -- $01222
          4643 => x"81", -- $01223
          4644 => x"81", -- $01224
          4645 => x"81", -- $01225
          4646 => x"81", -- $01226
          4647 => x"81", -- $01227
          4648 => x"81", -- $01228
          4649 => x"81", -- $01229
          4650 => x"81", -- $0122a
          4651 => x"81", -- $0122b
          4652 => x"81", -- $0122c
          4653 => x"81", -- $0122d
          4654 => x"81", -- $0122e
          4655 => x"81", -- $0122f
          4656 => x"81", -- $01230
          4657 => x"81", -- $01231
          4658 => x"81", -- $01232
          4659 => x"81", -- $01233
          4660 => x"81", -- $01234
          4661 => x"81", -- $01235
          4662 => x"81", -- $01236
          4663 => x"81", -- $01237
          4664 => x"81", -- $01238
          4665 => x"81", -- $01239
          4666 => x"81", -- $0123a
          4667 => x"80", -- $0123b
          4668 => x"80", -- $0123c
          4669 => x"80", -- $0123d
          4670 => x"80", -- $0123e
          4671 => x"81", -- $0123f
          4672 => x"81", -- $01240
          4673 => x"81", -- $01241
          4674 => x"80", -- $01242
          4675 => x"80", -- $01243
          4676 => x"80", -- $01244
          4677 => x"80", -- $01245
          4678 => x"80", -- $01246
          4679 => x"80", -- $01247
          4680 => x"80", -- $01248
          4681 => x"80", -- $01249
          4682 => x"80", -- $0124a
          4683 => x"80", -- $0124b
          4684 => x"80", -- $0124c
          4685 => x"80", -- $0124d
          4686 => x"80", -- $0124e
          4687 => x"80", -- $0124f
          4688 => x"80", -- $01250
          4689 => x"80", -- $01251
          4690 => x"80", -- $01252
          4691 => x"80", -- $01253
          4692 => x"80", -- $01254
          4693 => x"80", -- $01255
          4694 => x"80", -- $01256
          4695 => x"80", -- $01257
          4696 => x"80", -- $01258
          4697 => x"80", -- $01259
          4698 => x"80", -- $0125a
          4699 => x"80", -- $0125b
          4700 => x"80", -- $0125c
          4701 => x"80", -- $0125d
          4702 => x"80", -- $0125e
          4703 => x"80", -- $0125f
          4704 => x"80", -- $01260
          4705 => x"80", -- $01261
          4706 => x"80", -- $01262
          4707 => x"80", -- $01263
          4708 => x"80", -- $01264
          4709 => x"80", -- $01265
          4710 => x"80", -- $01266
          4711 => x"80", -- $01267
          4712 => x"80", -- $01268
          4713 => x"80", -- $01269
          4714 => x"80", -- $0126a
          4715 => x"80", -- $0126b
          4716 => x"80", -- $0126c
          4717 => x"80", -- $0126d
          4718 => x"80", -- $0126e
          4719 => x"80", -- $0126f
          4720 => x"80", -- $01270
          4721 => x"80", -- $01271
          4722 => x"80", -- $01272
          4723 => x"80", -- $01273
          4724 => x"80", -- $01274
          4725 => x"80", -- $01275
          4726 => x"80", -- $01276
          4727 => x"80", -- $01277
          4728 => x"80", -- $01278
          4729 => x"80", -- $01279
          4730 => x"80", -- $0127a
          4731 => x"80", -- $0127b
          4732 => x"80", -- $0127c
          4733 => x"80", -- $0127d
          4734 => x"80", -- $0127e
          4735 => x"80", -- $0127f
          4736 => x"80", -- $01280
          4737 => x"80", -- $01281
          4738 => x"80", -- $01282
          4739 => x"80", -- $01283
          4740 => x"80", -- $01284
          4741 => x"80", -- $01285
          4742 => x"80", -- $01286
          4743 => x"80", -- $01287
          4744 => x"80", -- $01288
          4745 => x"80", -- $01289
          4746 => x"80", -- $0128a
          4747 => x"80", -- $0128b
          4748 => x"80", -- $0128c
          4749 => x"80", -- $0128d
          4750 => x"80", -- $0128e
          4751 => x"80", -- $0128f
          4752 => x"80", -- $01290
          4753 => x"80", -- $01291
          4754 => x"80", -- $01292
          4755 => x"80", -- $01293
          4756 => x"80", -- $01294
          4757 => x"80", -- $01295
          4758 => x"80", -- $01296
          4759 => x"80", -- $01297
          4760 => x"80", -- $01298
          4761 => x"80", -- $01299
          4762 => x"80", -- $0129a
          4763 => x"80", -- $0129b
          4764 => x"80", -- $0129c
          4765 => x"80", -- $0129d
          4766 => x"80", -- $0129e
          4767 => x"80", -- $0129f
          4768 => x"80", -- $012a0
          4769 => x"80", -- $012a1
          4770 => x"7f", -- $012a2
          4771 => x"80", -- $012a3
          4772 => x"80", -- $012a4
          4773 => x"7f", -- $012a5
          4774 => x"7f", -- $012a6
          4775 => x"7f", -- $012a7
          4776 => x"7f", -- $012a8
          4777 => x"7f", -- $012a9
          4778 => x"7f", -- $012aa
          4779 => x"7f", -- $012ab
          4780 => x"7f", -- $012ac
          4781 => x"7f", -- $012ad
          4782 => x"7f", -- $012ae
          4783 => x"7f", -- $012af
          4784 => x"7f", -- $012b0
          4785 => x"7f", -- $012b1
          4786 => x"7f", -- $012b2
          4787 => x"7f", -- $012b3
          4788 => x"7f", -- $012b4
          4789 => x"7f", -- $012b5
          4790 => x"7f", -- $012b6
          4791 => x"7f", -- $012b7
          4792 => x"7e", -- $012b8
          4793 => x"7e", -- $012b9
          4794 => x"7e", -- $012ba
          4795 => x"7e", -- $012bb
          4796 => x"7e", -- $012bc
          4797 => x"7e", -- $012bd
          4798 => x"7e", -- $012be
          4799 => x"7e", -- $012bf
          4800 => x"7e", -- $012c0
          4801 => x"7e", -- $012c1
          4802 => x"7e", -- $012c2
          4803 => x"7e", -- $012c3
          4804 => x"7e", -- $012c4
          4805 => x"7e", -- $012c5
          4806 => x"7e", -- $012c6
          4807 => x"7e", -- $012c7
          4808 => x"7e", -- $012c8
          4809 => x"7e", -- $012c9
          4810 => x"7e", -- $012ca
          4811 => x"7e", -- $012cb
          4812 => x"7e", -- $012cc
          4813 => x"7e", -- $012cd
          4814 => x"7e", -- $012ce
          4815 => x"7e", -- $012cf
          4816 => x"7e", -- $012d0
          4817 => x"7e", -- $012d1
          4818 => x"7e", -- $012d2
          4819 => x"7e", -- $012d3
          4820 => x"7e", -- $012d4
          4821 => x"7e", -- $012d5
          4822 => x"7e", -- $012d6
          4823 => x"7e", -- $012d7
          4824 => x"7e", -- $012d8
          4825 => x"7e", -- $012d9
          4826 => x"7e", -- $012da
          4827 => x"7e", -- $012db
          4828 => x"7e", -- $012dc
          4829 => x"7e", -- $012dd
          4830 => x"7e", -- $012de
          4831 => x"7e", -- $012df
          4832 => x"7e", -- $012e0
          4833 => x"7e", -- $012e1
          4834 => x"7d", -- $012e2
          4835 => x"7d", -- $012e3
          4836 => x"7d", -- $012e4
          4837 => x"7d", -- $012e5
          4838 => x"7e", -- $012e6
          4839 => x"7e", -- $012e7
          4840 => x"7e", -- $012e8
          4841 => x"7e", -- $012e9
          4842 => x"7d", -- $012ea
          4843 => x"7d", -- $012eb
          4844 => x"7e", -- $012ec
          4845 => x"7e", -- $012ed
          4846 => x"7e", -- $012ee
          4847 => x"7e", -- $012ef
          4848 => x"7e", -- $012f0
          4849 => x"7d", -- $012f1
          4850 => x"7d", -- $012f2
          4851 => x"7e", -- $012f3
          4852 => x"7e", -- $012f4
          4853 => x"7e", -- $012f5
          4854 => x"7e", -- $012f6
          4855 => x"7e", -- $012f7
          4856 => x"7e", -- $012f8
          4857 => x"7e", -- $012f9
          4858 => x"7e", -- $012fa
          4859 => x"7e", -- $012fb
          4860 => x"7d", -- $012fc
          4861 => x"7e", -- $012fd
          4862 => x"7e", -- $012fe
          4863 => x"7e", -- $012ff
          4864 => x"7e", -- $01300
          4865 => x"7e", -- $01301
          4866 => x"7d", -- $01302
          4867 => x"7d", -- $01303
          4868 => x"7d", -- $01304
          4869 => x"7d", -- $01305
          4870 => x"7e", -- $01306
          4871 => x"7e", -- $01307
          4872 => x"7d", -- $01308
          4873 => x"7d", -- $01309
          4874 => x"7d", -- $0130a
          4875 => x"7d", -- $0130b
          4876 => x"7d", -- $0130c
          4877 => x"7d", -- $0130d
          4878 => x"7d", -- $0130e
          4879 => x"7d", -- $0130f
          4880 => x"7d", -- $01310
          4881 => x"7e", -- $01311
          4882 => x"7e", -- $01312
          4883 => x"7e", -- $01313
          4884 => x"7e", -- $01314
          4885 => x"7e", -- $01315
          4886 => x"7d", -- $01316
          4887 => x"7d", -- $01317
          4888 => x"7d", -- $01318
          4889 => x"7d", -- $01319
          4890 => x"7e", -- $0131a
          4891 => x"7e", -- $0131b
          4892 => x"7e", -- $0131c
          4893 => x"7e", -- $0131d
          4894 => x"7e", -- $0131e
          4895 => x"7e", -- $0131f
          4896 => x"7e", -- $01320
          4897 => x"7e", -- $01321
          4898 => x"7e", -- $01322
          4899 => x"7e", -- $01323
          4900 => x"7e", -- $01324
          4901 => x"7e", -- $01325
          4902 => x"7e", -- $01326
          4903 => x"7e", -- $01327
          4904 => x"7e", -- $01328
          4905 => x"7e", -- $01329
          4906 => x"7e", -- $0132a
          4907 => x"7e", -- $0132b
          4908 => x"7e", -- $0132c
          4909 => x"7e", -- $0132d
          4910 => x"7e", -- $0132e
          4911 => x"7e", -- $0132f
          4912 => x"7e", -- $01330
          4913 => x"7d", -- $01331
          4914 => x"7e", -- $01332
          4915 => x"7e", -- $01333
          4916 => x"7e", -- $01334
          4917 => x"7e", -- $01335
          4918 => x"7e", -- $01336
          4919 => x"7e", -- $01337
          4920 => x"7e", -- $01338
          4921 => x"7e", -- $01339
          4922 => x"7e", -- $0133a
          4923 => x"7e", -- $0133b
          4924 => x"7e", -- $0133c
          4925 => x"7e", -- $0133d
          4926 => x"7e", -- $0133e
          4927 => x"7e", -- $0133f
          4928 => x"7e", -- $01340
          4929 => x"7e", -- $01341
          4930 => x"7e", -- $01342
          4931 => x"7e", -- $01343
          4932 => x"7e", -- $01344
          4933 => x"7e", -- $01345
          4934 => x"7e", -- $01346
          4935 => x"7e", -- $01347
          4936 => x"7e", -- $01348
          4937 => x"7e", -- $01349
          4938 => x"7e", -- $0134a
          4939 => x"7e", -- $0134b
          4940 => x"7e", -- $0134c
          4941 => x"7e", -- $0134d
          4942 => x"7e", -- $0134e
          4943 => x"7e", -- $0134f
          4944 => x"7e", -- $01350
          4945 => x"7e", -- $01351
          4946 => x"7e", -- $01352
          4947 => x"7e", -- $01353
          4948 => x"7e", -- $01354
          4949 => x"7e", -- $01355
          4950 => x"7e", -- $01356
          4951 => x"7e", -- $01357
          4952 => x"7e", -- $01358
          4953 => x"7e", -- $01359
          4954 => x"7e", -- $0135a
          4955 => x"7e", -- $0135b
          4956 => x"7e", -- $0135c
          4957 => x"7e", -- $0135d
          4958 => x"7e", -- $0135e
          4959 => x"7e", -- $0135f
          4960 => x"7e", -- $01360
          4961 => x"7e", -- $01361
          4962 => x"7e", -- $01362
          4963 => x"7e", -- $01363
          4964 => x"7e", -- $01364
          4965 => x"7e", -- $01365
          4966 => x"7e", -- $01366
          4967 => x"7e", -- $01367
          4968 => x"7e", -- $01368
          4969 => x"7e", -- $01369
          4970 => x"7e", -- $0136a
          4971 => x"7e", -- $0136b
          4972 => x"7e", -- $0136c
          4973 => x"7e", -- $0136d
          4974 => x"7e", -- $0136e
          4975 => x"7e", -- $0136f
          4976 => x"7e", -- $01370
          4977 => x"7e", -- $01371
          4978 => x"7e", -- $01372
          4979 => x"7e", -- $01373
          4980 => x"7e", -- $01374
          4981 => x"7e", -- $01375
          4982 => x"7e", -- $01376
          4983 => x"7e", -- $01377
          4984 => x"7e", -- $01378
          4985 => x"7e", -- $01379
          4986 => x"7e", -- $0137a
          4987 => x"7e", -- $0137b
          4988 => x"7e", -- $0137c
          4989 => x"7e", -- $0137d
          4990 => x"7e", -- $0137e
          4991 => x"7e", -- $0137f
          4992 => x"7e", -- $01380
          4993 => x"7e", -- $01381
          4994 => x"7e", -- $01382
          4995 => x"7e", -- $01383
          4996 => x"7e", -- $01384
          4997 => x"7e", -- $01385
          4998 => x"7e", -- $01386
          4999 => x"7e", -- $01387
          5000 => x"7e", -- $01388
          5001 => x"7e", -- $01389
          5002 => x"7e", -- $0138a
          5003 => x"7e", -- $0138b
          5004 => x"7e", -- $0138c
          5005 => x"7e", -- $0138d
          5006 => x"7e", -- $0138e
          5007 => x"7e", -- $0138f
          5008 => x"7e", -- $01390
          5009 => x"7e", -- $01391
          5010 => x"7e", -- $01392
          5011 => x"7e", -- $01393
          5012 => x"7e", -- $01394
          5013 => x"7e", -- $01395
          5014 => x"7e", -- $01396
          5015 => x"7e", -- $01397
          5016 => x"7e", -- $01398
          5017 => x"7e", -- $01399
          5018 => x"7e", -- $0139a
          5019 => x"7e", -- $0139b
          5020 => x"7e", -- $0139c
          5021 => x"7e", -- $0139d
          5022 => x"7e", -- $0139e
          5023 => x"7e", -- $0139f
          5024 => x"7e", -- $013a0
          5025 => x"7e", -- $013a1
          5026 => x"7e", -- $013a2
          5027 => x"7e", -- $013a3
          5028 => x"7e", -- $013a4
          5029 => x"7e", -- $013a5
          5030 => x"7e", -- $013a6
          5031 => x"7e", -- $013a7
          5032 => x"7e", -- $013a8
          5033 => x"7e", -- $013a9
          5034 => x"7e", -- $013aa
          5035 => x"7e", -- $013ab
          5036 => x"7e", -- $013ac
          5037 => x"7e", -- $013ad
          5038 => x"7e", -- $013ae
          5039 => x"7e", -- $013af
          5040 => x"7f", -- $013b0
          5041 => x"7f", -- $013b1
          5042 => x"7f", -- $013b2
          5043 => x"7e", -- $013b3
          5044 => x"7f", -- $013b4
          5045 => x"7f", -- $013b5
          5046 => x"7f", -- $013b6
          5047 => x"7e", -- $013b7
          5048 => x"7f", -- $013b8
          5049 => x"7f", -- $013b9
          5050 => x"7f", -- $013ba
          5051 => x"7e", -- $013bb
          5052 => x"7e", -- $013bc
          5053 => x"7e", -- $013bd
          5054 => x"7d", -- $013be
          5055 => x"7e", -- $013bf
          5056 => x"7d", -- $013c0
          5057 => x"7e", -- $013c1
          5058 => x"7d", -- $013c2
          5059 => x"7d", -- $013c3
          5060 => x"7d", -- $013c4
          5061 => x"7c", -- $013c5
          5062 => x"7d", -- $013c6
          5063 => x"7c", -- $013c7
          5064 => x"7d", -- $013c8
          5065 => x"7d", -- $013c9
          5066 => x"7e", -- $013ca
          5067 => x"7d", -- $013cb
          5068 => x"7e", -- $013cc
          5069 => x"7f", -- $013cd
          5070 => x"7f", -- $013ce
          5071 => x"80", -- $013cf
          5072 => x"80", -- $013d0
          5073 => x"80", -- $013d1
          5074 => x"80", -- $013d2
          5075 => x"82", -- $013d3
          5076 => x"82", -- $013d4
          5077 => x"82", -- $013d5
          5078 => x"83", -- $013d6
          5079 => x"83", -- $013d7
          5080 => x"83", -- $013d8
          5081 => x"83", -- $013d9
          5082 => x"82", -- $013da
          5083 => x"82", -- $013db
          5084 => x"81", -- $013dc
          5085 => x"80", -- $013dd
          5086 => x"80", -- $013de
          5087 => x"7f", -- $013df
          5088 => x"80", -- $013e0
          5089 => x"7e", -- $013e1
          5090 => x"7f", -- $013e2
          5091 => x"7e", -- $013e3
          5092 => x"7e", -- $013e4
          5093 => x"7e", -- $013e5
          5094 => x"7e", -- $013e6
          5095 => x"7f", -- $013e7
          5096 => x"7e", -- $013e8
          5097 => x"80", -- $013e9
          5098 => x"80", -- $013ea
          5099 => x"80", -- $013eb
          5100 => x"80", -- $013ec
          5101 => x"80", -- $013ed
          5102 => x"81", -- $013ee
          5103 => x"82", -- $013ef
          5104 => x"82", -- $013f0
          5105 => x"82", -- $013f1
          5106 => x"82", -- $013f2
          5107 => x"82", -- $013f3
          5108 => x"82", -- $013f4
          5109 => x"82", -- $013f5
          5110 => x"81", -- $013f6
          5111 => x"81", -- $013f7
          5112 => x"81", -- $013f8
          5113 => x"80", -- $013f9
          5114 => x"80", -- $013fa
          5115 => x"80", -- $013fb
          5116 => x"80", -- $013fc
          5117 => x"80", -- $013fd
          5118 => x"7f", -- $013fe
          5119 => x"7f", -- $013ff
          5120 => x"7f", -- $01400
          5121 => x"7e", -- $01401
          5122 => x"7e", -- $01402
          5123 => x"7e", -- $01403
          5124 => x"7e", -- $01404
          5125 => x"7e", -- $01405
          5126 => x"7e", -- $01406
          5127 => x"7e", -- $01407
          5128 => x"7f", -- $01408
          5129 => x"7f", -- $01409
          5130 => x"80", -- $0140a
          5131 => x"80", -- $0140b
          5132 => x"81", -- $0140c
          5133 => x"82", -- $0140d
          5134 => x"82", -- $0140e
          5135 => x"84", -- $0140f
          5136 => x"85", -- $01410
          5137 => x"86", -- $01411
          5138 => x"86", -- $01412
          5139 => x"87", -- $01413
          5140 => x"88", -- $01414
          5141 => x"88", -- $01415
          5142 => x"88", -- $01416
          5143 => x"88", -- $01417
          5144 => x"88", -- $01418
          5145 => x"87", -- $01419
          5146 => x"87", -- $0141a
          5147 => x"86", -- $0141b
          5148 => x"85", -- $0141c
          5149 => x"83", -- $0141d
          5150 => x"82", -- $0141e
          5151 => x"81", -- $0141f
          5152 => x"80", -- $01420
          5153 => x"7f", -- $01421
          5154 => x"7e", -- $01422
          5155 => x"7e", -- $01423
          5156 => x"7d", -- $01424
          5157 => x"7c", -- $01425
          5158 => x"7c", -- $01426
          5159 => x"7c", -- $01427
          5160 => x"7c", -- $01428
          5161 => x"7c", -- $01429
          5162 => x"7d", -- $0142a
          5163 => x"7d", -- $0142b
          5164 => x"7d", -- $0142c
          5165 => x"7e", -- $0142d
          5166 => x"7e", -- $0142e
          5167 => x"7f", -- $0142f
          5168 => x"80", -- $01430
          5169 => x"80", -- $01431
          5170 => x"80", -- $01432
          5171 => x"81", -- $01433
          5172 => x"81", -- $01434
          5173 => x"81", -- $01435
          5174 => x"82", -- $01436
          5175 => x"82", -- $01437
          5176 => x"82", -- $01438
          5177 => x"82", -- $01439
          5178 => x"83", -- $0143a
          5179 => x"83", -- $0143b
          5180 => x"83", -- $0143c
          5181 => x"83", -- $0143d
          5182 => x"84", -- $0143e
          5183 => x"84", -- $0143f
          5184 => x"84", -- $01440
          5185 => x"85", -- $01441
          5186 => x"85", -- $01442
          5187 => x"86", -- $01443
          5188 => x"86", -- $01444
          5189 => x"87", -- $01445
          5190 => x"87", -- $01446
          5191 => x"88", -- $01447
          5192 => x"88", -- $01448
          5193 => x"87", -- $01449
          5194 => x"88", -- $0144a
          5195 => x"86", -- $0144b
          5196 => x"86", -- $0144c
          5197 => x"85", -- $0144d
          5198 => x"84", -- $0144e
          5199 => x"84", -- $0144f
          5200 => x"82", -- $01450
          5201 => x"81", -- $01451
          5202 => x"80", -- $01452
          5203 => x"80", -- $01453
          5204 => x"80", -- $01454
          5205 => x"7f", -- $01455
          5206 => x"7f", -- $01456
          5207 => x"7f", -- $01457
          5208 => x"7f", -- $01458
          5209 => x"7e", -- $01459
          5210 => x"7f", -- $0145a
          5211 => x"7e", -- $0145b
          5212 => x"7e", -- $0145c
          5213 => x"7e", -- $0145d
          5214 => x"7e", -- $0145e
          5215 => x"7e", -- $0145f
          5216 => x"7d", -- $01460
          5217 => x"7f", -- $01461
          5218 => x"7f", -- $01462
          5219 => x"80", -- $01463
          5220 => x"80", -- $01464
          5221 => x"80", -- $01465
          5222 => x"81", -- $01466
          5223 => x"81", -- $01467
          5224 => x"82", -- $01468
          5225 => x"81", -- $01469
          5226 => x"82", -- $0146a
          5227 => x"82", -- $0146b
          5228 => x"82", -- $0146c
          5229 => x"82", -- $0146d
          5230 => x"82", -- $0146e
          5231 => x"82", -- $0146f
          5232 => x"81", -- $01470
          5233 => x"82", -- $01471
          5234 => x"81", -- $01472
          5235 => x"81", -- $01473
          5236 => x"82", -- $01474
          5237 => x"82", -- $01475
          5238 => x"83", -- $01476
          5239 => x"83", -- $01477
          5240 => x"85", -- $01478
          5241 => x"84", -- $01479
          5242 => x"86", -- $0147a
          5243 => x"86", -- $0147b
          5244 => x"87", -- $0147c
          5245 => x"88", -- $0147d
          5246 => x"87", -- $0147e
          5247 => x"87", -- $0147f
          5248 => x"87", -- $01480
          5249 => x"87", -- $01481
          5250 => x"86", -- $01482
          5251 => x"87", -- $01483
          5252 => x"85", -- $01484
          5253 => x"86", -- $01485
          5254 => x"84", -- $01486
          5255 => x"83", -- $01487
          5256 => x"84", -- $01488
          5257 => x"83", -- $01489
          5258 => x"83", -- $0148a
          5259 => x"82", -- $0148b
          5260 => x"81", -- $0148c
          5261 => x"81", -- $0148d
          5262 => x"80", -- $0148e
          5263 => x"80", -- $0148f
          5264 => x"80", -- $01490
          5265 => x"7f", -- $01491
          5266 => x"7e", -- $01492
          5267 => x"7e", -- $01493
          5268 => x"7d", -- $01494
          5269 => x"7d", -- $01495
          5270 => x"7d", -- $01496
          5271 => x"7d", -- $01497
          5272 => x"7e", -- $01498
          5273 => x"7e", -- $01499
          5274 => x"7f", -- $0149a
          5275 => x"80", -- $0149b
          5276 => x"80", -- $0149c
          5277 => x"81", -- $0149d
          5278 => x"81", -- $0149e
          5279 => x"82", -- $0149f
          5280 => x"82", -- $014a0
          5281 => x"82", -- $014a1
          5282 => x"82", -- $014a2
          5283 => x"82", -- $014a3
          5284 => x"81", -- $014a4
          5285 => x"81", -- $014a5
          5286 => x"80", -- $014a6
          5287 => x"80", -- $014a7
          5288 => x"80", -- $014a8
          5289 => x"80", -- $014a9
          5290 => x"80", -- $014aa
          5291 => x"80", -- $014ab
          5292 => x"80", -- $014ac
          5293 => x"81", -- $014ad
          5294 => x"82", -- $014ae
          5295 => x"83", -- $014af
          5296 => x"84", -- $014b0
          5297 => x"85", -- $014b1
          5298 => x"87", -- $014b2
          5299 => x"87", -- $014b3
          5300 => x"88", -- $014b4
          5301 => x"89", -- $014b5
          5302 => x"89", -- $014b6
          5303 => x"8b", -- $014b7
          5304 => x"8a", -- $014b8
          5305 => x"8b", -- $014b9
          5306 => x"8a", -- $014ba
          5307 => x"8a", -- $014bb
          5308 => x"8a", -- $014bc
          5309 => x"89", -- $014bd
          5310 => x"8a", -- $014be
          5311 => x"88", -- $014bf
          5312 => x"88", -- $014c0
          5313 => x"86", -- $014c1
          5314 => x"85", -- $014c2
          5315 => x"83", -- $014c3
          5316 => x"81", -- $014c4
          5317 => x"81", -- $014c5
          5318 => x"7f", -- $014c6
          5319 => x"7f", -- $014c7
          5320 => x"7d", -- $014c8
          5321 => x"7d", -- $014c9
          5322 => x"7c", -- $014ca
          5323 => x"7b", -- $014cb
          5324 => x"7b", -- $014cc
          5325 => x"7b", -- $014cd
          5326 => x"7c", -- $014ce
          5327 => x"7d", -- $014cf
          5328 => x"7d", -- $014d0
          5329 => x"7f", -- $014d1
          5330 => x"80", -- $014d2
          5331 => x"80", -- $014d3
          5332 => x"82", -- $014d4
          5333 => x"83", -- $014d5
          5334 => x"84", -- $014d6
          5335 => x"84", -- $014d7
          5336 => x"85", -- $014d8
          5337 => x"85", -- $014d9
          5338 => x"85", -- $014da
          5339 => x"84", -- $014db
          5340 => x"84", -- $014dc
          5341 => x"84", -- $014dd
          5342 => x"82", -- $014de
          5343 => x"83", -- $014df
          5344 => x"82", -- $014e0
          5345 => x"82", -- $014e1
          5346 => x"81", -- $014e2
          5347 => x"81", -- $014e3
          5348 => x"82", -- $014e4
          5349 => x"81", -- $014e5
          5350 => x"82", -- $014e6
          5351 => x"82", -- $014e7
          5352 => x"82", -- $014e8
          5353 => x"84", -- $014e9
          5354 => x"82", -- $014ea
          5355 => x"84", -- $014eb
          5356 => x"83", -- $014ec
          5357 => x"85", -- $014ed
          5358 => x"86", -- $014ee
          5359 => x"86", -- $014ef
          5360 => x"87", -- $014f0
          5361 => x"87", -- $014f1
          5362 => x"89", -- $014f2
          5363 => x"87", -- $014f3
          5364 => x"8a", -- $014f4
          5365 => x"87", -- $014f5
          5366 => x"8b", -- $014f6
          5367 => x"89", -- $014f7
          5368 => x"88", -- $014f8
          5369 => x"8b", -- $014f9
          5370 => x"86", -- $014fa
          5371 => x"88", -- $014fb
          5372 => x"85", -- $014fc
          5373 => x"86", -- $014fd
          5374 => x"84", -- $014fe
          5375 => x"83", -- $014ff
          5376 => x"82", -- $01500
          5377 => x"81", -- $01501
          5378 => x"80", -- $01502
          5379 => x"7e", -- $01503
          5380 => x"80", -- $01504
          5381 => x"7d", -- $01505
          5382 => x"7e", -- $01506
          5383 => x"7d", -- $01507
          5384 => x"7c", -- $01508
          5385 => x"7f", -- $01509
          5386 => x"7c", -- $0150a
          5387 => x"80", -- $0150b
          5388 => x"7f", -- $0150c
          5389 => x"81", -- $0150d
          5390 => x"81", -- $0150e
          5391 => x"81", -- $0150f
          5392 => x"84", -- $01510
          5393 => x"81", -- $01511
          5394 => x"84", -- $01512
          5395 => x"81", -- $01513
          5396 => x"83", -- $01514
          5397 => x"81", -- $01515
          5398 => x"80", -- $01516
          5399 => x"82", -- $01517
          5400 => x"7f", -- $01518
          5401 => x"81", -- $01519
          5402 => x"7e", -- $0151a
          5403 => x"80", -- $0151b
          5404 => x"7f", -- $0151c
          5405 => x"7d", -- $0151d
          5406 => x"7f", -- $0151e
          5407 => x"7d", -- $0151f
          5408 => x"80", -- $01520
          5409 => x"7e", -- $01521
          5410 => x"80", -- $01522
          5411 => x"80", -- $01523
          5412 => x"80", -- $01524
          5413 => x"82", -- $01525
          5414 => x"82", -- $01526
          5415 => x"85", -- $01527
          5416 => x"85", -- $01528
          5417 => x"85", -- $01529
          5418 => x"85", -- $0152a
          5419 => x"89", -- $0152b
          5420 => x"88", -- $0152c
          5421 => x"87", -- $0152d
          5422 => x"8b", -- $0152e
          5423 => x"87", -- $0152f
          5424 => x"8d", -- $01530
          5425 => x"87", -- $01531
          5426 => x"89", -- $01532
          5427 => x"8c", -- $01533
          5428 => x"86", -- $01534
          5429 => x"89", -- $01535
          5430 => x"85", -- $01536
          5431 => x"86", -- $01537
          5432 => x"83", -- $01538
          5433 => x"82", -- $01539
          5434 => x"81", -- $0153a
          5435 => x"80", -- $0153b
          5436 => x"7e", -- $0153c
          5437 => x"7c", -- $0153d
          5438 => x"7e", -- $0153e
          5439 => x"7a", -- $0153f
          5440 => x"7a", -- $01540
          5441 => x"78", -- $01541
          5442 => x"7a", -- $01542
          5443 => x"7a", -- $01543
          5444 => x"78", -- $01544
          5445 => x"7c", -- $01545
          5446 => x"7c", -- $01546
          5447 => x"7e", -- $01547
          5448 => x"7d", -- $01548
          5449 => x"80", -- $01549
          5450 => x"80", -- $0154a
          5451 => x"80", -- $0154b
          5452 => x"81", -- $0154c
          5453 => x"80", -- $0154d
          5454 => x"82", -- $0154e
          5455 => x"80", -- $0154f
          5456 => x"81", -- $01550
          5457 => x"80", -- $01551
          5458 => x"80", -- $01552
          5459 => x"7f", -- $01553
          5460 => x"7e", -- $01554
          5461 => x"7f", -- $01555
          5462 => x"7d", -- $01556
          5463 => x"7d", -- $01557
          5464 => x"7d", -- $01558
          5465 => x"7c", -- $01559
          5466 => x"7c", -- $0155a
          5467 => x"7c", -- $0155b
          5468 => x"7d", -- $0155c
          5469 => x"7d", -- $0155d
          5470 => x"7d", -- $0155e
          5471 => x"7d", -- $0155f
          5472 => x"7e", -- $01560
          5473 => x"7f", -- $01561
          5474 => x"7f", -- $01562
          5475 => x"81", -- $01563
          5476 => x"82", -- $01564
          5477 => x"82", -- $01565
          5478 => x"81", -- $01566
          5479 => x"86", -- $01567
          5480 => x"86", -- $01568
          5481 => x"84", -- $01569
          5482 => x"8a", -- $0156a
          5483 => x"85", -- $0156b
          5484 => x"8c", -- $0156c
          5485 => x"88", -- $0156d
          5486 => x"87", -- $0156e
          5487 => x"8e", -- $0156f
          5488 => x"86", -- $01570
          5489 => x"89", -- $01571
          5490 => x"87", -- $01572
          5491 => x"86", -- $01573
          5492 => x"86", -- $01574
          5493 => x"82", -- $01575
          5494 => x"81", -- $01576
          5495 => x"82", -- $01577
          5496 => x"7f", -- $01578
          5497 => x"7c", -- $01579
          5498 => x"7e", -- $0157a
          5499 => x"79", -- $0157b
          5500 => x"7a", -- $0157c
          5501 => x"78", -- $0157d
          5502 => x"78", -- $0157e
          5503 => x"79", -- $0157f
          5504 => x"77", -- $01580
          5505 => x"7a", -- $01581
          5506 => x"7b", -- $01582
          5507 => x"7c", -- $01583
          5508 => x"7c", -- $01584
          5509 => x"7e", -- $01585
          5510 => x"7f", -- $01586
          5511 => x"7f", -- $01587
          5512 => x"7e", -- $01588
          5513 => x"7f", -- $01589
          5514 => x"80", -- $0158a
          5515 => x"7d", -- $0158b
          5516 => x"7e", -- $0158c
          5517 => x"7e", -- $0158d
          5518 => x"7c", -- $0158e
          5519 => x"7c", -- $0158f
          5520 => x"7b", -- $01590
          5521 => x"7c", -- $01591
          5522 => x"7a", -- $01592
          5523 => x"7a", -- $01593
          5524 => x"7b", -- $01594
          5525 => x"7b", -- $01595
          5526 => x"7b", -- $01596
          5527 => x"7b", -- $01597
          5528 => x"7d", -- $01598
          5529 => x"7d", -- $01599
          5530 => x"7d", -- $0159a
          5531 => x"7e", -- $0159b
          5532 => x"7f", -- $0159c
          5533 => x"80", -- $0159d
          5534 => x"80", -- $0159e
          5535 => x"82", -- $0159f
          5536 => x"83", -- $015a0
          5537 => x"84", -- $015a1
          5538 => x"86", -- $015a2
          5539 => x"84", -- $015a3
          5540 => x"86", -- $015a4
          5541 => x"8b", -- $015a5
          5542 => x"85", -- $015a6
          5543 => x"89", -- $015a7
          5544 => x"8b", -- $015a8
          5545 => x"88", -- $015a9
          5546 => x"8d", -- $015aa
          5547 => x"86", -- $015ab
          5548 => x"89", -- $015ac
          5549 => x"8c", -- $015ad
          5550 => x"83", -- $015ae
          5551 => x"86", -- $015af
          5552 => x"86", -- $015b0
          5553 => x"80", -- $015b1
          5554 => x"81", -- $015b2
          5555 => x"80", -- $015b3
          5556 => x"7d", -- $015b4
          5557 => x"80", -- $015b5
          5558 => x"79", -- $015b6
          5559 => x"7a", -- $015b7
          5560 => x"7c", -- $015b8
          5561 => x"75", -- $015b9
          5562 => x"77", -- $015ba
          5563 => x"77", -- $015bb
          5564 => x"77", -- $015bc
          5565 => x"78", -- $015bd
          5566 => x"77", -- $015be
          5567 => x"79", -- $015bf
          5568 => x"7c", -- $015c0
          5569 => x"7a", -- $015c1
          5570 => x"7c", -- $015c2
          5571 => x"7f", -- $015c3
          5572 => x"7d", -- $015c4
          5573 => x"7e", -- $015c5
          5574 => x"7e", -- $015c6
          5575 => x"7e", -- $015c7
          5576 => x"7e", -- $015c8
          5577 => x"7b", -- $015c9
          5578 => x"7c", -- $015ca
          5579 => x"7d", -- $015cb
          5580 => x"7a", -- $015cc
          5581 => x"7a", -- $015cd
          5582 => x"7a", -- $015ce
          5583 => x"79", -- $015cf
          5584 => x"78", -- $015d0
          5585 => x"78", -- $015d1
          5586 => x"79", -- $015d2
          5587 => x"79", -- $015d3
          5588 => x"79", -- $015d4
          5589 => x"7a", -- $015d5
          5590 => x"7c", -- $015d6
          5591 => x"7c", -- $015d7
          5592 => x"7c", -- $015d8
          5593 => x"7e", -- $015d9
          5594 => x"7f", -- $015da
          5595 => x"80", -- $015db
          5596 => x"80", -- $015dc
          5597 => x"82", -- $015dd
          5598 => x"83", -- $015de
          5599 => x"84", -- $015df
          5600 => x"85", -- $015e0
          5601 => x"85", -- $015e1
          5602 => x"87", -- $015e2
          5603 => x"8b", -- $015e3
          5604 => x"86", -- $015e4
          5605 => x"8a", -- $015e5
          5606 => x"8c", -- $015e6
          5607 => x"87", -- $015e7
          5608 => x"8b", -- $015e8
          5609 => x"88", -- $015e9
          5610 => x"88", -- $015ea
          5611 => x"8b", -- $015eb
          5612 => x"84", -- $015ec
          5613 => x"84", -- $015ed
          5614 => x"87", -- $015ee
          5615 => x"80", -- $015ef
          5616 => x"80", -- $015f0
          5617 => x"81", -- $015f1
          5618 => x"7c", -- $015f2
          5619 => x"7c", -- $015f3
          5620 => x"7a", -- $015f4
          5621 => x"77", -- $015f5
          5622 => x"79", -- $015f6
          5623 => x"75", -- $015f7
          5624 => x"73", -- $015f8
          5625 => x"76", -- $015f9
          5626 => x"75", -- $015fa
          5627 => x"73", -- $015fb
          5628 => x"77", -- $015fc
          5629 => x"77", -- $015fd
          5630 => x"78", -- $015fe
          5631 => x"79", -- $015ff
          5632 => x"7a", -- $01600
          5633 => x"7c", -- $01601
          5634 => x"7a", -- $01602
          5635 => x"7b", -- $01603
          5636 => x"7c", -- $01604
          5637 => x"7c", -- $01605
          5638 => x"7b", -- $01606
          5639 => x"7a", -- $01607
          5640 => x"7b", -- $01608
          5641 => x"79", -- $01609
          5642 => x"78", -- $0160a
          5643 => x"78", -- $0160b
          5644 => x"78", -- $0160c
          5645 => x"77", -- $0160d
          5646 => x"77", -- $0160e
          5647 => x"78", -- $0160f
          5648 => x"78", -- $01610
          5649 => x"79", -- $01611
          5650 => x"79", -- $01612
          5651 => x"7a", -- $01613
          5652 => x"7c", -- $01614
          5653 => x"7c", -- $01615
          5654 => x"7d", -- $01616
          5655 => x"7f", -- $01617
          5656 => x"80", -- $01618
          5657 => x"80", -- $01619
          5658 => x"81", -- $0161a
          5659 => x"83", -- $0161b
          5660 => x"83", -- $0161c
          5661 => x"85", -- $0161d
          5662 => x"86", -- $0161e
          5663 => x"88", -- $0161f
          5664 => x"87", -- $01620
          5665 => x"85", -- $01621
          5666 => x"8c", -- $01622
          5667 => x"8a", -- $01623
          5668 => x"86", -- $01624
          5669 => x"8a", -- $01625
          5670 => x"8b", -- $01626
          5671 => x"88", -- $01627
          5672 => x"86", -- $01628
          5673 => x"86", -- $01629
          5674 => x"88", -- $0162a
          5675 => x"84", -- $0162b
          5676 => x"80", -- $0162c
          5677 => x"82", -- $0162d
          5678 => x"81", -- $0162e
          5679 => x"7d", -- $0162f
          5680 => x"7b", -- $01630
          5681 => x"7b", -- $01631
          5682 => x"7a", -- $01632
          5683 => x"76", -- $01633
          5684 => x"75", -- $01634
          5685 => x"76", -- $01635
          5686 => x"75", -- $01636
          5687 => x"74", -- $01637
          5688 => x"73", -- $01638
          5689 => x"76", -- $01639
          5690 => x"77", -- $0163a
          5691 => x"75", -- $0163b
          5692 => x"77", -- $0163c
          5693 => x"7a", -- $0163d
          5694 => x"7b", -- $0163e
          5695 => x"78", -- $0163f
          5696 => x"7c", -- $01640
          5697 => x"7d", -- $01641
          5698 => x"7b", -- $01642
          5699 => x"7a", -- $01643
          5700 => x"7b", -- $01644
          5701 => x"7b", -- $01645
          5702 => x"78", -- $01646
          5703 => x"77", -- $01647
          5704 => x"77", -- $01648
          5705 => x"76", -- $01649
          5706 => x"75", -- $0164a
          5707 => x"73", -- $0164b
          5708 => x"74", -- $0164c
          5709 => x"75", -- $0164d
          5710 => x"74", -- $0164e
          5711 => x"74", -- $0164f
          5712 => x"77", -- $01650
          5713 => x"79", -- $01651
          5714 => x"79", -- $01652
          5715 => x"7a", -- $01653
          5716 => x"7d", -- $01654
          5717 => x"80", -- $01655
          5718 => x"7f", -- $01656
          5719 => x"80", -- $01657
          5720 => x"84", -- $01658
          5721 => x"84", -- $01659
          5722 => x"84", -- $0165a
          5723 => x"85", -- $0165b
          5724 => x"89", -- $0165c
          5725 => x"89", -- $0165d
          5726 => x"88", -- $0165e
          5727 => x"8b", -- $0165f
          5728 => x"8c", -- $01660
          5729 => x"89", -- $01661
          5730 => x"89", -- $01662
          5731 => x"8d", -- $01663
          5732 => x"8b", -- $01664
          5733 => x"88", -- $01665
          5734 => x"88", -- $01666
          5735 => x"8b", -- $01667
          5736 => x"88", -- $01668
          5737 => x"82", -- $01669
          5738 => x"84", -- $0166a
          5739 => x"85", -- $0166b
          5740 => x"80", -- $0166c
          5741 => x"7d", -- $0166d
          5742 => x"7e", -- $0166e
          5743 => x"7e", -- $0166f
          5744 => x"79", -- $01670
          5745 => x"77", -- $01671
          5746 => x"76", -- $01672
          5747 => x"76", -- $01673
          5748 => x"74", -- $01674
          5749 => x"72", -- $01675
          5750 => x"73", -- $01676
          5751 => x"74", -- $01677
          5752 => x"73", -- $01678
          5753 => x"73", -- $01679
          5754 => x"76", -- $0167a
          5755 => x"77", -- $0167b
          5756 => x"77", -- $0167c
          5757 => x"79", -- $0167d
          5758 => x"7b", -- $0167e
          5759 => x"7d", -- $0167f
          5760 => x"7b", -- $01680
          5761 => x"7d", -- $01681
          5762 => x"7d", -- $01682
          5763 => x"7c", -- $01683
          5764 => x"7a", -- $01684
          5765 => x"79", -- $01685
          5766 => x"7a", -- $01686
          5767 => x"77", -- $01687
          5768 => x"76", -- $01688
          5769 => x"74", -- $01689
          5770 => x"75", -- $0168a
          5771 => x"74", -- $0168b
          5772 => x"72", -- $0168c
          5773 => x"74", -- $0168d
          5774 => x"76", -- $0168e
          5775 => x"77", -- $0168f
          5776 => x"78", -- $01690
          5777 => x"7a", -- $01691
          5778 => x"7d", -- $01692
          5779 => x"7f", -- $01693
          5780 => x"80", -- $01694
          5781 => x"82", -- $01695
          5782 => x"84", -- $01696
          5783 => x"87", -- $01697
          5784 => x"88", -- $01698
          5785 => x"89", -- $01699
          5786 => x"8a", -- $0169a
          5787 => x"8d", -- $0169b
          5788 => x"8d", -- $0169c
          5789 => x"8c", -- $0169d
          5790 => x"8d", -- $0169e
          5791 => x"8e", -- $0169f
          5792 => x"8f", -- $016a0
          5793 => x"8d", -- $016a1
          5794 => x"8a", -- $016a2
          5795 => x"89", -- $016a3
          5796 => x"8d", -- $016a4
          5797 => x"8c", -- $016a5
          5798 => x"87", -- $016a6
          5799 => x"85", -- $016a7
          5800 => x"89", -- $016a8
          5801 => x"89", -- $016a9
          5802 => x"83", -- $016aa
          5803 => x"80", -- $016ab
          5804 => x"82", -- $016ac
          5805 => x"82", -- $016ad
          5806 => x"7e", -- $016ae
          5807 => x"7a", -- $016af
          5808 => x"7a", -- $016b0
          5809 => x"7a", -- $016b1
          5810 => x"78", -- $016b2
          5811 => x"75", -- $016b3
          5812 => x"74", -- $016b4
          5813 => x"74", -- $016b5
          5814 => x"75", -- $016b6
          5815 => x"75", -- $016b7
          5816 => x"74", -- $016b8
          5817 => x"74", -- $016b9
          5818 => x"78", -- $016ba
          5819 => x"7b", -- $016bb
          5820 => x"7a", -- $016bc
          5821 => x"7a", -- $016bd
          5822 => x"7e", -- $016be
          5823 => x"80", -- $016bf
          5824 => x"7f", -- $016c0
          5825 => x"7d", -- $016c1
          5826 => x"7e", -- $016c2
          5827 => x"7e", -- $016c3
          5828 => x"7c", -- $016c4
          5829 => x"7a", -- $016c5
          5830 => x"78", -- $016c6
          5831 => x"76", -- $016c7
          5832 => x"75", -- $016c8
          5833 => x"75", -- $016c9
          5834 => x"73", -- $016ca
          5835 => x"72", -- $016cb
          5836 => x"73", -- $016cc
          5837 => x"76", -- $016cd
          5838 => x"77", -- $016ce
          5839 => x"79", -- $016cf
          5840 => x"7c", -- $016d0
          5841 => x"80", -- $016d1
          5842 => x"82", -- $016d2
          5843 => x"85", -- $016d3
          5844 => x"87", -- $016d4
          5845 => x"8a", -- $016d5
          5846 => x"8c", -- $016d6
          5847 => x"8e", -- $016d7
          5848 => x"90", -- $016d8
          5849 => x"8f", -- $016d9
          5850 => x"8f", -- $016da
          5851 => x"8f", -- $016db
          5852 => x"90", -- $016dc
          5853 => x"8d", -- $016dd
          5854 => x"8c", -- $016de
          5855 => x"8d", -- $016df
          5856 => x"8e", -- $016e0
          5857 => x"8c", -- $016e1
          5858 => x"88", -- $016e2
          5859 => x"86", -- $016e3
          5860 => x"88", -- $016e4
          5861 => x"88", -- $016e5
          5862 => x"89", -- $016e6
          5863 => x"87", -- $016e7
          5864 => x"85", -- $016e8
          5865 => x"85", -- $016e9
          5866 => x"86", -- $016ea
          5867 => x"85", -- $016eb
          5868 => x"82", -- $016ec
          5869 => x"80", -- $016ed
          5870 => x"7f", -- $016ee
          5871 => x"7e", -- $016ef
          5872 => x"7c", -- $016f0
          5873 => x"79", -- $016f1
          5874 => x"76", -- $016f2
          5875 => x"74", -- $016f3
          5876 => x"74", -- $016f4
          5877 => x"74", -- $016f5
          5878 => x"75", -- $016f6
          5879 => x"75", -- $016f7
          5880 => x"74", -- $016f8
          5881 => x"76", -- $016f9
          5882 => x"78", -- $016fa
          5883 => x"7c", -- $016fb
          5884 => x"7e", -- $016fc
          5885 => x"7e", -- $016fd
          5886 => x"7e", -- $016fe
          5887 => x"80", -- $016ff
          5888 => x"81", -- $01700
          5889 => x"80", -- $01701
          5890 => x"7f", -- $01702
          5891 => x"7c", -- $01703
          5892 => x"7b", -- $01704
          5893 => x"7a", -- $01705
          5894 => x"78", -- $01706
          5895 => x"75", -- $01707
          5896 => x"71", -- $01708
          5897 => x"70", -- $01709
          5898 => x"71", -- $0170a
          5899 => x"72", -- $0170b
          5900 => x"73", -- $0170c
          5901 => x"74", -- $0170d
          5902 => x"77", -- $0170e
          5903 => x"7a", -- $0170f
          5904 => x"7f", -- $01710
          5905 => x"83", -- $01711
          5906 => x"86", -- $01712
          5907 => x"88", -- $01713
          5908 => x"8b", -- $01714
          5909 => x"8e", -- $01715
          5910 => x"90", -- $01716
          5911 => x"92", -- $01717
          5912 => x"91", -- $01718
          5913 => x"90", -- $01719
          5914 => x"8e", -- $0171a
          5915 => x"8d", -- $0171b
          5916 => x"8d", -- $0171c
          5917 => x"8b", -- $0171d
          5918 => x"88", -- $0171e
          5919 => x"86", -- $0171f
          5920 => x"88", -- $01720
          5921 => x"89", -- $01721
          5922 => x"8a", -- $01722
          5923 => x"8a", -- $01723
          5924 => x"88", -- $01724
          5925 => x"88", -- $01725
          5926 => x"88", -- $01726
          5927 => x"8a", -- $01727
          5928 => x"8c", -- $01728
          5929 => x"8a", -- $01729
          5930 => x"89", -- $0172a
          5931 => x"86", -- $0172b
          5932 => x"85", -- $0172c
          5933 => x"83", -- $0172d
          5934 => x"82", -- $0172e
          5935 => x"7f", -- $0172f
          5936 => x"7b", -- $01730
          5937 => x"77", -- $01731
          5938 => x"74", -- $01732
          5939 => x"73", -- $01733
          5940 => x"72", -- $01734
          5941 => x"72", -- $01735
          5942 => x"71", -- $01736
          5943 => x"72", -- $01737
          5944 => x"74", -- $01738
          5945 => x"77", -- $01739
          5946 => x"7a", -- $0173a
          5947 => x"7d", -- $0173b
          5948 => x"7f", -- $0173c
          5949 => x"80", -- $0173d
          5950 => x"82", -- $0173e
          5951 => x"84", -- $0173f
          5952 => x"84", -- $01740
          5953 => x"84", -- $01741
          5954 => x"82", -- $01742
          5955 => x"80", -- $01743
          5956 => x"7d", -- $01744
          5957 => x"7b", -- $01745
          5958 => x"78", -- $01746
          5959 => x"75", -- $01747
          5960 => x"72", -- $01748
          5961 => x"6f", -- $01749
          5962 => x"6f", -- $0174a
          5963 => x"6e", -- $0174b
          5964 => x"70", -- $0174c
          5965 => x"75", -- $0174d
          5966 => x"78", -- $0174e
          5967 => x"7c", -- $0174f
          5968 => x"80", -- $01750
          5969 => x"85", -- $01751
          5970 => x"8a", -- $01752
          5971 => x"8f", -- $01753
          5972 => x"93", -- $01754
          5973 => x"94", -- $01755
          5974 => x"95", -- $01756
          5975 => x"94", -- $01757
          5976 => x"92", -- $01758
          5977 => x"91", -- $01759
          5978 => x"8e", -- $0175a
          5979 => x"8c", -- $0175b
          5980 => x"88", -- $0175c
          5981 => x"85", -- $0175d
          5982 => x"84", -- $0175e
          5983 => x"83", -- $0175f
          5984 => x"83", -- $01760
          5985 => x"83", -- $01761
          5986 => x"85", -- $01762
          5987 => x"88", -- $01763
          5988 => x"8c", -- $01764
          5989 => x"8f", -- $01765
          5990 => x"91", -- $01766
          5991 => x"94", -- $01767
          5992 => x"93", -- $01768
          5993 => x"91", -- $01769
          5994 => x"8e", -- $0176a
          5995 => x"8c", -- $0176b
          5996 => x"8a", -- $0176c
          5997 => x"87", -- $0176d
          5998 => x"84", -- $0176e
          5999 => x"81", -- $0176f
          6000 => x"7d", -- $01770
          6001 => x"79", -- $01771
          6002 => x"77", -- $01772
          6003 => x"76", -- $01773
          6004 => x"75", -- $01774
          6005 => x"75", -- $01775
          6006 => x"75", -- $01776
          6007 => x"76", -- $01777
          6008 => x"76", -- $01778
          6009 => x"78", -- $01779
          6010 => x"7b", -- $0177a
          6011 => x"7e", -- $0177b
          6012 => x"80", -- $0177c
          6013 => x"82", -- $0177d
          6014 => x"83", -- $0177e
          6015 => x"82", -- $0177f
          6016 => x"82", -- $01780
          6017 => x"81", -- $01781
          6018 => x"82", -- $01782
          6019 => x"81", -- $01783
          6020 => x"80", -- $01784
          6021 => x"7f", -- $01785
          6022 => x"7b", -- $01786
          6023 => x"79", -- $01787
          6024 => x"76", -- $01788
          6025 => x"75", -- $01789
          6026 => x"75", -- $0178a
          6027 => x"75", -- $0178b
          6028 => x"75", -- $0178c
          6029 => x"76", -- $0178d
          6030 => x"78", -- $0178e
          6031 => x"7a", -- $0178f
          6032 => x"7f", -- $01790
          6033 => x"83", -- $01791
          6034 => x"87", -- $01792
          6035 => x"8c", -- $01793
          6036 => x"8f", -- $01794
          6037 => x"91", -- $01795
          6038 => x"93", -- $01796
          6039 => x"93", -- $01797
          6040 => x"93", -- $01798
          6041 => x"92", -- $01799
          6042 => x"90", -- $0179a
          6043 => x"8d", -- $0179b
          6044 => x"89", -- $0179c
          6045 => x"85", -- $0179d
          6046 => x"83", -- $0179e
          6047 => x"81", -- $0179f
          6048 => x"80", -- $017a0
          6049 => x"80", -- $017a1
          6050 => x"80", -- $017a2
          6051 => x"83", -- $017a3
          6052 => x"86", -- $017a4
          6053 => x"89", -- $017a5
          6054 => x"8c", -- $017a6
          6055 => x"8e", -- $017a7
          6056 => x"90", -- $017a8
          6057 => x"91", -- $017a9
          6058 => x"92", -- $017aa
          6059 => x"91", -- $017ab
          6060 => x"90", -- $017ac
          6061 => x"8c", -- $017ad
          6062 => x"87", -- $017ae
          6063 => x"82", -- $017af
          6064 => x"7d", -- $017b0
          6065 => x"7b", -- $017b1
          6066 => x"79", -- $017b2
          6067 => x"7a", -- $017b3
          6068 => x"7a", -- $017b4
          6069 => x"7a", -- $017b5
          6070 => x"7b", -- $017b6
          6071 => x"7a", -- $017b7
          6072 => x"7a", -- $017b8
          6073 => x"7a", -- $017b9
          6074 => x"7c", -- $017ba
          6075 => x"7e", -- $017bb
          6076 => x"7f", -- $017bc
          6077 => x"7f", -- $017bd
          6078 => x"7e", -- $017be
          6079 => x"7c", -- $017bf
          6080 => x"7b", -- $017c0
          6081 => x"7c", -- $017c1
          6082 => x"7d", -- $017c2
          6083 => x"7f", -- $017c3
          6084 => x"80", -- $017c4
          6085 => x"80", -- $017c5
          6086 => x"80", -- $017c6
          6087 => x"7f", -- $017c7
          6088 => x"7f", -- $017c8
          6089 => x"7f", -- $017c9
          6090 => x"80", -- $017ca
          6091 => x"80", -- $017cb
          6092 => x"80", -- $017cc
          6093 => x"80", -- $017cd
          6094 => x"7d", -- $017ce
          6095 => x"7b", -- $017cf
          6096 => x"7a", -- $017d0
          6097 => x"7a", -- $017d1
          6098 => x"7b", -- $017d2
          6099 => x"7d", -- $017d3
          6100 => x"80", -- $017d4
          6101 => x"82", -- $017d5
          6102 => x"85", -- $017d6
          6103 => x"87", -- $017d7
          6104 => x"8a", -- $017d8
          6105 => x"8c", -- $017d9
          6106 => x"8f", -- $017da
          6107 => x"90", -- $017db
          6108 => x"90", -- $017dc
          6109 => x"8f", -- $017dd
          6110 => x"8c", -- $017de
          6111 => x"89", -- $017df
          6112 => x"86", -- $017e0
          6113 => x"83", -- $017e1
          6114 => x"81", -- $017e2
          6115 => x"80", -- $017e3
          6116 => x"80", -- $017e4
          6117 => x"80", -- $017e5
          6118 => x"80", -- $017e6
          6119 => x"81", -- $017e7
          6120 => x"83", -- $017e8
          6121 => x"85", -- $017e9
          6122 => x"87", -- $017ea
          6123 => x"8a", -- $017eb
          6124 => x"8b", -- $017ec
          6125 => x"8c", -- $017ed
          6126 => x"8c", -- $017ee
          6127 => x"8a", -- $017ef
          6128 => x"88", -- $017f0
          6129 => x"86", -- $017f1
          6130 => x"83", -- $017f2
          6131 => x"81", -- $017f3
          6132 => x"80", -- $017f4
          6133 => x"7f", -- $017f5
          6134 => x"7d", -- $017f6
          6135 => x"7c", -- $017f7
          6136 => x"7b", -- $017f8
          6137 => x"7b", -- $017f9
          6138 => x"7c", -- $017fa
          6139 => x"7f", -- $017fb
          6140 => x"81", -- $017fc
          6141 => x"83", -- $017fd
          6142 => x"85", -- $017fe
          6143 => x"84", -- $017ff
          6144 => x"81", -- $01800
          6145 => x"7f", -- $01801
          6146 => x"7c", -- $01802
          6147 => x"7a", -- $01803
          6148 => x"78", -- $01804
          6149 => x"78", -- $01805
          6150 => x"78", -- $01806
          6151 => x"78", -- $01807
          6152 => x"79", -- $01808
          6153 => x"7a", -- $01809
          6154 => x"7d", -- $0180a
          6155 => x"80", -- $0180b
          6156 => x"82", -- $0180c
          6157 => x"85", -- $0180d
          6158 => x"88", -- $0180e
          6159 => x"88", -- $0180f
          6160 => x"89", -- $01810
          6161 => x"88", -- $01811
          6162 => x"86", -- $01812
          6163 => x"83", -- $01813
          6164 => x"80", -- $01814
          6165 => x"7f", -- $01815
          6166 => x"7d", -- $01816
          6167 => x"7c", -- $01817
          6168 => x"7a", -- $01818
          6169 => x"7b", -- $01819
          6170 => x"7c", -- $0181a
          6171 => x"7e", -- $0181b
          6172 => x"80", -- $0181c
          6173 => x"84", -- $0181d
          6174 => x"87", -- $0181e
          6175 => x"8a", -- $0181f
          6176 => x"8c", -- $01820
          6177 => x"8d", -- $01821
          6178 => x"8d", -- $01822
          6179 => x"8b", -- $01823
          6180 => x"89", -- $01824
          6181 => x"85", -- $01825
          6182 => x"81", -- $01826
          6183 => x"7f", -- $01827
          6184 => x"7c", -- $01828
          6185 => x"7b", -- $01829
          6186 => x"7b", -- $0182a
          6187 => x"7c", -- $0182b
          6188 => x"7d", -- $0182c
          6189 => x"7f", -- $0182d
          6190 => x"81", -- $0182e
          6191 => x"83", -- $0182f
          6192 => x"86", -- $01830
          6193 => x"87", -- $01831
          6194 => x"89", -- $01832
          6195 => x"89", -- $01833
          6196 => x"88", -- $01834
          6197 => x"88", -- $01835
          6198 => x"85", -- $01836
          6199 => x"83", -- $01837
          6200 => x"80", -- $01838
          6201 => x"80", -- $01839
          6202 => x"7e", -- $0183a
          6203 => x"7d", -- $0183b
          6204 => x"7d", -- $0183c
          6205 => x"7e", -- $0183d
          6206 => x"80", -- $0183e
          6207 => x"80", -- $0183f
          6208 => x"81", -- $01840
          6209 => x"82", -- $01841
          6210 => x"82", -- $01842
          6211 => x"82", -- $01843
          6212 => x"82", -- $01844
          6213 => x"82", -- $01845
          6214 => x"82", -- $01846
          6215 => x"82", -- $01847
          6216 => x"81", -- $01848
          6217 => x"81", -- $01849
          6218 => x"80", -- $0184a
          6219 => x"7d", -- $0184b
          6220 => x"7b", -- $0184c
          6221 => x"7a", -- $0184d
          6222 => x"79", -- $0184e
          6223 => x"7a", -- $0184f
          6224 => x"7c", -- $01850
          6225 => x"7e", -- $01851
          6226 => x"80", -- $01852
          6227 => x"83", -- $01853
          6228 => x"85", -- $01854
          6229 => x"86", -- $01855
          6230 => x"86", -- $01856
          6231 => x"86", -- $01857
          6232 => x"86", -- $01858
          6233 => x"85", -- $01859
          6234 => x"84", -- $0185a
          6235 => x"82", -- $0185b
          6236 => x"80", -- $0185c
          6237 => x"7f", -- $0185d
          6238 => x"7d", -- $0185e
          6239 => x"7c", -- $0185f
          6240 => x"7b", -- $01860
          6241 => x"7b", -- $01861
          6242 => x"7c", -- $01862
          6243 => x"7d", -- $01863
          6244 => x"7e", -- $01864
          6245 => x"7f", -- $01865
          6246 => x"80", -- $01866
          6247 => x"81", -- $01867
          6248 => x"82", -- $01868
          6249 => x"82", -- $01869
          6250 => x"82", -- $0186a
          6251 => x"82", -- $0186b
          6252 => x"82", -- $0186c
          6253 => x"80", -- $0186d
          6254 => x"80", -- $0186e
          6255 => x"7e", -- $0186f
          6256 => x"7d", -- $01870
          6257 => x"7b", -- $01871
          6258 => x"7b", -- $01872
          6259 => x"7b", -- $01873
          6260 => x"7c", -- $01874
          6261 => x"7d", -- $01875
          6262 => x"7f", -- $01876
          6263 => x"80", -- $01877
          6264 => x"83", -- $01878
          6265 => x"84", -- $01879
          6266 => x"85", -- $0187a
          6267 => x"86", -- $0187b
          6268 => x"85", -- $0187c
          6269 => x"84", -- $0187d
          6270 => x"83", -- $0187e
          6271 => x"82", -- $0187f
          6272 => x"81", -- $01880
          6273 => x"80", -- $01881
          6274 => x"80", -- $01882
          6275 => x"7f", -- $01883
          6276 => x"7e", -- $01884
          6277 => x"7f", -- $01885
          6278 => x"80", -- $01886
          6279 => x"81", -- $01887
          6280 => x"83", -- $01888
          6281 => x"85", -- $01889
          6282 => x"85", -- $0188a
          6283 => x"85", -- $0188b
          6284 => x"83", -- $0188c
          6285 => x"81", -- $0188d
          6286 => x"80", -- $0188e
          6287 => x"7f", -- $0188f
          6288 => x"80", -- $01890
          6289 => x"80", -- $01891
          6290 => x"81", -- $01892
          6291 => x"82", -- $01893
          6292 => x"81", -- $01894
          6293 => x"80", -- $01895
          6294 => x"7f", -- $01896
          6295 => x"7d", -- $01897
          6296 => x"7b", -- $01898
          6297 => x"7b", -- $01899
          6298 => x"7c", -- $0189a
          6299 => x"7d", -- $0189b
          6300 => x"7f", -- $0189c
          6301 => x"80", -- $0189d
          6302 => x"81", -- $0189e
          6303 => x"80", -- $0189f
          6304 => x"80", -- $018a0
          6305 => x"7f", -- $018a1
          6306 => x"7d", -- $018a2
          6307 => x"7c", -- $018a3
          6308 => x"7c", -- $018a4
          6309 => x"7c", -- $018a5
          6310 => x"7d", -- $018a6
          6311 => x"7d", -- $018a7
          6312 => x"7d", -- $018a8
          6313 => x"7d", -- $018a9
          6314 => x"7d", -- $018aa
          6315 => x"7c", -- $018ab
          6316 => x"7b", -- $018ac
          6317 => x"7c", -- $018ad
          6318 => x"7b", -- $018ae
          6319 => x"7d", -- $018af
          6320 => x"7e", -- $018b0
          6321 => x"7e", -- $018b1
          6322 => x"7f", -- $018b2
          6323 => x"7e", -- $018b3
          6324 => x"7d", -- $018b4
          6325 => x"7c", -- $018b5
          6326 => x"7b", -- $018b6
          6327 => x"7b", -- $018b7
          6328 => x"7b", -- $018b8
          6329 => x"7c", -- $018b9
          6330 => x"7d", -- $018ba
          6331 => x"7e", -- $018bb
          6332 => x"7e", -- $018bc
          6333 => x"7e", -- $018bd
          6334 => x"7e", -- $018be
          6335 => x"7f", -- $018bf
          6336 => x"80", -- $018c0
          6337 => x"80", -- $018c1
          6338 => x"81", -- $018c2
          6339 => x"82", -- $018c3
          6340 => x"83", -- $018c4
          6341 => x"83", -- $018c5
          6342 => x"82", -- $018c6
          6343 => x"81", -- $018c7
          6344 => x"80", -- $018c8
          6345 => x"7f", -- $018c9
          6346 => x"7e", -- $018ca
          6347 => x"7f", -- $018cb
          6348 => x"7e", -- $018cc
          6349 => x"7f", -- $018cd
          6350 => x"80", -- $018ce
          6351 => x"80", -- $018cf
          6352 => x"81", -- $018d0
          6353 => x"82", -- $018d1
          6354 => x"83", -- $018d2
          6355 => x"84", -- $018d3
          6356 => x"85", -- $018d4
          6357 => x"85", -- $018d5
          6358 => x"85", -- $018d6
          6359 => x"84", -- $018d7
          6360 => x"82", -- $018d8
          6361 => x"7f", -- $018d9
          6362 => x"7d", -- $018da
          6363 => x"7b", -- $018db
          6364 => x"79", -- $018dc
          6365 => x"7a", -- $018dd
          6366 => x"7b", -- $018de
          6367 => x"7d", -- $018df
          6368 => x"7f", -- $018e0
          6369 => x"80", -- $018e1
          6370 => x"80", -- $018e2
          6371 => x"7e", -- $018e3
          6372 => x"7d", -- $018e4
          6373 => x"7b", -- $018e5
          6374 => x"7a", -- $018e6
          6375 => x"79", -- $018e7
          6376 => x"79", -- $018e8
          6377 => x"7a", -- $018e9
          6378 => x"7b", -- $018ea
          6379 => x"7c", -- $018eb
          6380 => x"7c", -- $018ec
          6381 => x"7c", -- $018ed
          6382 => x"7b", -- $018ee
          6383 => x"7a", -- $018ef
          6384 => x"7a", -- $018f0
          6385 => x"7a", -- $018f1
          6386 => x"7b", -- $018f2
          6387 => x"7d", -- $018f3
          6388 => x"7e", -- $018f4
          6389 => x"7f", -- $018f5
          6390 => x"7f", -- $018f6
          6391 => x"7e", -- $018f7
          6392 => x"7d", -- $018f8
          6393 => x"7b", -- $018f9
          6394 => x"79", -- $018fa
          6395 => x"79", -- $018fb
          6396 => x"79", -- $018fc
          6397 => x"7a", -- $018fd
          6398 => x"7c", -- $018fe
          6399 => x"7d", -- $018ff
          6400 => x"7e", -- $01900
          6401 => x"7f", -- $01901
          6402 => x"80", -- $01902
          6403 => x"80", -- $01903
          6404 => x"80", -- $01904
          6405 => x"80", -- $01905
          6406 => x"81", -- $01906
          6407 => x"81", -- $01907
          6408 => x"81", -- $01908
          6409 => x"81", -- $01909
          6410 => x"80", -- $0190a
          6411 => x"80", -- $0190b
          6412 => x"7f", -- $0190c
          6413 => x"7e", -- $0190d
          6414 => x"7e", -- $0190e
          6415 => x"7e", -- $0190f
          6416 => x"7f", -- $01910
          6417 => x"80", -- $01911
          6418 => x"81", -- $01912
          6419 => x"82", -- $01913
          6420 => x"84", -- $01914
          6421 => x"84", -- $01915
          6422 => x"84", -- $01916
          6423 => x"83", -- $01917
          6424 => x"82", -- $01918
          6425 => x"81", -- $01919
          6426 => x"81", -- $0191a
          6427 => x"80", -- $0191b
          6428 => x"80", -- $0191c
          6429 => x"80", -- $0191d
          6430 => x"80", -- $0191e
          6431 => x"81", -- $0191f
          6432 => x"81", -- $01920
          6433 => x"81", -- $01921
          6434 => x"80", -- $01922
          6435 => x"80", -- $01923
          6436 => x"7e", -- $01924
          6437 => x"7e", -- $01925
          6438 => x"7d", -- $01926
          6439 => x"7e", -- $01927
          6440 => x"7f", -- $01928
          6441 => x"80", -- $01929
          6442 => x"81", -- $0192a
          6443 => x"81", -- $0192b
          6444 => x"80", -- $0192c
          6445 => x"7e", -- $0192d
          6446 => x"7b", -- $0192e
          6447 => x"78", -- $0192f
          6448 => x"75", -- $01930
          6449 => x"74", -- $01931
          6450 => x"74", -- $01932
          6451 => x"75", -- $01933
          6452 => x"77", -- $01934
          6453 => x"7b", -- $01935
          6454 => x"7d", -- $01936
          6455 => x"7f", -- $01937
          6456 => x"80", -- $01938
          6457 => x"80", -- $01939
          6458 => x"80", -- $0193a
          6459 => x"80", -- $0193b
          6460 => x"7f", -- $0193c
          6461 => x"7f", -- $0193d
          6462 => x"7f", -- $0193e
          6463 => x"7f", -- $0193f
          6464 => x"7f", -- $01940
          6465 => x"7d", -- $01941
          6466 => x"7d", -- $01942
          6467 => x"7b", -- $01943
          6468 => x"7b", -- $01944
          6469 => x"7a", -- $01945
          6470 => x"7b", -- $01946
          6471 => x"7c", -- $01947
          6472 => x"7e", -- $01948
          6473 => x"80", -- $01949
          6474 => x"81", -- $0194a
          6475 => x"83", -- $0194b
          6476 => x"83", -- $0194c
          6477 => x"83", -- $0194d
          6478 => x"82", -- $0194e
          6479 => x"80", -- $0194f
          6480 => x"80", -- $01950
          6481 => x"7e", -- $01951
          6482 => x"7d", -- $01952
          6483 => x"7c", -- $01953
          6484 => x"7d", -- $01954
          6485 => x"7d", -- $01955
          6486 => x"7d", -- $01956
          6487 => x"7e", -- $01957
          6488 => x"7e", -- $01958
          6489 => x"7f", -- $01959
          6490 => x"80", -- $0195a
          6491 => x"81", -- $0195b
          6492 => x"81", -- $0195c
          6493 => x"82", -- $0195d
          6494 => x"82", -- $0195e
          6495 => x"81", -- $0195f
          6496 => x"81", -- $01960
          6497 => x"80", -- $01961
          6498 => x"7f", -- $01962
          6499 => x"7e", -- $01963
          6500 => x"7d", -- $01964
          6501 => x"7d", -- $01965
          6502 => x"7d", -- $01966
          6503 => x"7e", -- $01967
          6504 => x"7f", -- $01968
          6505 => x"80", -- $01969
          6506 => x"82", -- $0196a
          6507 => x"83", -- $0196b
          6508 => x"85", -- $0196c
          6509 => x"84", -- $0196d
          6510 => x"84", -- $0196e
          6511 => x"82", -- $0196f
          6512 => x"80", -- $01970
          6513 => x"7f", -- $01971
          6514 => x"7c", -- $01972
          6515 => x"7c", -- $01973
          6516 => x"7c", -- $01974
          6517 => x"7d", -- $01975
          6518 => x"7e", -- $01976
          6519 => x"7e", -- $01977
          6520 => x"7e", -- $01978
          6521 => x"7d", -- $01979
          6522 => x"7c", -- $0197a
          6523 => x"79", -- $0197b
          6524 => x"78", -- $0197c
          6525 => x"77", -- $0197d
          6526 => x"77", -- $0197e
          6527 => x"78", -- $0197f
          6528 => x"7a", -- $01980
          6529 => x"7d", -- $01981
          6530 => x"7f", -- $01982
          6531 => x"80", -- $01983
          6532 => x"80", -- $01984
          6533 => x"80", -- $01985
          6534 => x"80", -- $01986
          6535 => x"7f", -- $01987
          6536 => x"7e", -- $01988
          6537 => x"7e", -- $01989
          6538 => x"7e", -- $0198a
          6539 => x"7e", -- $0198b
          6540 => x"7e", -- $0198c
          6541 => x"7e", -- $0198d
          6542 => x"7e", -- $0198e
          6543 => x"7e", -- $0198f
          6544 => x"7d", -- $01990
          6545 => x"7d", -- $01991
          6546 => x"7d", -- $01992
          6547 => x"7d", -- $01993
          6548 => x"7e", -- $01994
          6549 => x"7f", -- $01995
          6550 => x"7f", -- $01996
          6551 => x"80", -- $01997
          6552 => x"80", -- $01998
          6553 => x"80", -- $01999
          6554 => x"80", -- $0199a
          6555 => x"80", -- $0199b
          6556 => x"80", -- $0199c
          6557 => x"7f", -- $0199d
          6558 => x"7e", -- $0199e
          6559 => x"7d", -- $0199f
          6560 => x"7d", -- $019a0
          6561 => x"7c", -- $019a1
          6562 => x"7d", -- $019a2
          6563 => x"7d", -- $019a3
          6564 => x"7e", -- $019a4
          6565 => x"7f", -- $019a5
          6566 => x"80", -- $019a6
          6567 => x"80", -- $019a7
          6568 => x"81", -- $019a8
          6569 => x"81", -- $019a9
          6570 => x"81", -- $019aa
          6571 => x"81", -- $019ab
          6572 => x"80", -- $019ac
          6573 => x"80", -- $019ad
          6574 => x"7f", -- $019ae
          6575 => x"7e", -- $019af
          6576 => x"7e", -- $019b0
          6577 => x"7f", -- $019b1
          6578 => x"7f", -- $019b2
          6579 => x"80", -- $019b3
          6580 => x"80", -- $019b4
          6581 => x"81", -- $019b5
          6582 => x"81", -- $019b6
          6583 => x"82", -- $019b7
          6584 => x"82", -- $019b8
          6585 => x"82", -- $019b9
          6586 => x"83", -- $019ba
          6587 => x"83", -- $019bb
          6588 => x"84", -- $019bc
          6589 => x"84", -- $019bd
          6590 => x"84", -- $019be
          6591 => x"83", -- $019bf
          6592 => x"81", -- $019c0
          6593 => x"80", -- $019c1
          6594 => x"7f", -- $019c2
          6595 => x"7e", -- $019c3
          6596 => x"7e", -- $019c4
          6597 => x"7f", -- $019c5
          6598 => x"80", -- $019c6
          6599 => x"80", -- $019c7
          6600 => x"81", -- $019c8
          6601 => x"80", -- $019c9
          6602 => x"80", -- $019ca
          6603 => x"7e", -- $019cb
          6604 => x"7b", -- $019cc
          6605 => x"78", -- $019cd
          6606 => x"76", -- $019ce
          6607 => x"76", -- $019cf
          6608 => x"77", -- $019d0
          6609 => x"79", -- $019d1
          6610 => x"7c", -- $019d2
          6611 => x"7f", -- $019d3
          6612 => x"81", -- $019d4
          6613 => x"82", -- $019d5
          6614 => x"83", -- $019d6
          6615 => x"83", -- $019d7
          6616 => x"83", -- $019d8
          6617 => x"82", -- $019d9
          6618 => x"82", -- $019da
          6619 => x"82", -- $019db
          6620 => x"81", -- $019dc
          6621 => x"80", -- $019dd
          6622 => x"80", -- $019de
          6623 => x"7e", -- $019df
          6624 => x"7c", -- $019e0
          6625 => x"7a", -- $019e1
          6626 => x"79", -- $019e2
          6627 => x"79", -- $019e3
          6628 => x"7a", -- $019e4
          6629 => x"7c", -- $019e5
          6630 => x"7e", -- $019e6
          6631 => x"80", -- $019e7
          6632 => x"82", -- $019e8
          6633 => x"84", -- $019e9
          6634 => x"84", -- $019ea
          6635 => x"84", -- $019eb
          6636 => x"82", -- $019ec
          6637 => x"80", -- $019ed
          6638 => x"80", -- $019ee
          6639 => x"7e", -- $019ef
          6640 => x"7d", -- $019f0
          6641 => x"7d", -- $019f1
          6642 => x"7d", -- $019f2
          6643 => x"7d", -- $019f3
          6644 => x"7e", -- $019f4
          6645 => x"7f", -- $019f5
          6646 => x"80", -- $019f6
          6647 => x"81", -- $019f7
          6648 => x"83", -- $019f8
          6649 => x"84", -- $019f9
          6650 => x"85", -- $019fa
          6651 => x"85", -- $019fb
          6652 => x"84", -- $019fc
          6653 => x"83", -- $019fd
          6654 => x"82", -- $019fe
          6655 => x"81", -- $019ff
          6656 => x"80", -- $01a00
          6657 => x"80", -- $01a01
          6658 => x"81", -- $01a02
          6659 => x"82", -- $01a03
          6660 => x"83", -- $01a04
          6661 => x"84", -- $01a05
          6662 => x"85", -- $01a06
          6663 => x"85", -- $01a07
          6664 => x"85", -- $01a08
          6665 => x"85", -- $01a09
          6666 => x"84", -- $01a0a
          6667 => x"83", -- $01a0b
          6668 => x"83", -- $01a0c
          6669 => x"83", -- $01a0d
          6670 => x"83", -- $01a0e
          6671 => x"83", -- $01a0f
          6672 => x"83", -- $01a10
          6673 => x"82", -- $01a11
          6674 => x"80", -- $01a12
          6675 => x"7f", -- $01a13
          6676 => x"7c", -- $01a14
          6677 => x"79", -- $01a15
          6678 => x"77", -- $01a16
          6679 => x"75", -- $01a17
          6680 => x"75", -- $01a18
          6681 => x"76", -- $01a19
          6682 => x"79", -- $01a1a
          6683 => x"7c", -- $01a1b
          6684 => x"7f", -- $01a1c
          6685 => x"82", -- $01a1d
          6686 => x"84", -- $01a1e
          6687 => x"85", -- $01a1f
          6688 => x"85", -- $01a20
          6689 => x"85", -- $01a21
          6690 => x"83", -- $01a22
          6691 => x"81", -- $01a23
          6692 => x"80", -- $01a24
          6693 => x"7e", -- $01a25
          6694 => x"7d", -- $01a26
          6695 => x"7c", -- $01a27
          6696 => x"7c", -- $01a28
          6697 => x"7b", -- $01a29
          6698 => x"7c", -- $01a2a
          6699 => x"7d", -- $01a2b
          6700 => x"7e", -- $01a2c
          6701 => x"7f", -- $01a2d
          6702 => x"80", -- $01a2e
          6703 => x"81", -- $01a2f
          6704 => x"82", -- $01a30
          6705 => x"83", -- $01a31
          6706 => x"84", -- $01a32
          6707 => x"84", -- $01a33
          6708 => x"83", -- $01a34
          6709 => x"82", -- $01a35
          6710 => x"81", -- $01a36
          6711 => x"80", -- $01a37
          6712 => x"7e", -- $01a38
          6713 => x"7d", -- $01a39
          6714 => x"7c", -- $01a3a
          6715 => x"7c", -- $01a3b
          6716 => x"7d", -- $01a3c
          6717 => x"7f", -- $01a3d
          6718 => x"80", -- $01a3e
          6719 => x"82", -- $01a3f
          6720 => x"84", -- $01a40
          6721 => x"86", -- $01a41
          6722 => x"87", -- $01a42
          6723 => x"88", -- $01a43
          6724 => x"87", -- $01a44
          6725 => x"86", -- $01a45
          6726 => x"84", -- $01a46
          6727 => x"82", -- $01a47
          6728 => x"80", -- $01a48
          6729 => x"7e", -- $01a49
          6730 => x"7d", -- $01a4a
          6731 => x"7d", -- $01a4b
          6732 => x"7d", -- $01a4c
          6733 => x"7f", -- $01a4d
          6734 => x"81", -- $01a4e
          6735 => x"84", -- $01a4f
          6736 => x"86", -- $01a50
          6737 => x"88", -- $01a51
          6738 => x"89", -- $01a52
          6739 => x"89", -- $01a53
          6740 => x"88", -- $01a54
          6741 => x"87", -- $01a55
          6742 => x"86", -- $01a56
          6743 => x"85", -- $01a57
          6744 => x"85", -- $01a58
          6745 => x"84", -- $01a59
          6746 => x"82", -- $01a5a
          6747 => x"81", -- $01a5b
          6748 => x"80", -- $01a5c
          6749 => x"7f", -- $01a5d
          6750 => x"7f", -- $01a5e
          6751 => x"7f", -- $01a5f
          6752 => x"80", -- $01a60
          6753 => x"81", -- $01a61
          6754 => x"82", -- $01a62
          6755 => x"83", -- $01a63
          6756 => x"82", -- $01a64
          6757 => x"80", -- $01a65
          6758 => x"7e", -- $01a66
          6759 => x"7b", -- $01a67
          6760 => x"77", -- $01a68
          6761 => x"75", -- $01a69
          6762 => x"75", -- $01a6a
          6763 => x"76", -- $01a6b
          6764 => x"79", -- $01a6c
          6765 => x"7c", -- $01a6d
          6766 => x"80", -- $01a6e
          6767 => x"84", -- $01a6f
          6768 => x"86", -- $01a70
          6769 => x"88", -- $01a71
          6770 => x"88", -- $01a72
          6771 => x"88", -- $01a73
          6772 => x"86", -- $01a74
          6773 => x"85", -- $01a75
          6774 => x"84", -- $01a76
          6775 => x"83", -- $01a77
          6776 => x"82", -- $01a78
          6777 => x"80", -- $01a79
          6778 => x"7f", -- $01a7a
          6779 => x"7c", -- $01a7b
          6780 => x"7b", -- $01a7c
          6781 => x"7a", -- $01a7d
          6782 => x"7a", -- $01a7e
          6783 => x"7d", -- $01a7f
          6784 => x"7f", -- $01a80
          6785 => x"81", -- $01a81
          6786 => x"84", -- $01a82
          6787 => x"86", -- $01a83
          6788 => x"87", -- $01a84
          6789 => x"87", -- $01a85
          6790 => x"87", -- $01a86
          6791 => x"85", -- $01a87
          6792 => x"84", -- $01a88
          6793 => x"82", -- $01a89
          6794 => x"80", -- $01a8a
          6795 => x"80", -- $01a8b
          6796 => x"7f", -- $01a8c
          6797 => x"7f", -- $01a8d
          6798 => x"7f", -- $01a8e
          6799 => x"80", -- $01a8f
          6800 => x"81", -- $01a90
          6801 => x"82", -- $01a91
          6802 => x"84", -- $01a92
          6803 => x"85", -- $01a93
          6804 => x"86", -- $01a94
          6805 => x"86", -- $01a95
          6806 => x"86", -- $01a96
          6807 => x"85", -- $01a97
          6808 => x"84", -- $01a98
          6809 => x"83", -- $01a99
          6810 => x"81", -- $01a9a
          6811 => x"81", -- $01a9b
          6812 => x"81", -- $01a9c
          6813 => x"82", -- $01a9d
          6814 => x"84", -- $01a9e
          6815 => x"85", -- $01a9f
          6816 => x"87", -- $01aa0
          6817 => x"88", -- $01aa1
          6818 => x"89", -- $01aa2
          6819 => x"88", -- $01aa3
          6820 => x"87", -- $01aa4
          6821 => x"86", -- $01aa5
          6822 => x"84", -- $01aa6
          6823 => x"83", -- $01aa7
          6824 => x"82", -- $01aa8
          6825 => x"82", -- $01aa9
          6826 => x"82", -- $01aaa
          6827 => x"83", -- $01aab
          6828 => x"84", -- $01aac
          6829 => x"83", -- $01aad
          6830 => x"82", -- $01aae
          6831 => x"80", -- $01aaf
          6832 => x"7d", -- $01ab0
          6833 => x"7a", -- $01ab1
          6834 => x"77", -- $01ab2
          6835 => x"77", -- $01ab3
          6836 => x"77", -- $01ab4
          6837 => x"79", -- $01ab5
          6838 => x"7c", -- $01ab6
          6839 => x"7f", -- $01ab7
          6840 => x"81", -- $01ab8
          6841 => x"84", -- $01ab9
          6842 => x"85", -- $01aba
          6843 => x"85", -- $01abb
          6844 => x"85", -- $01abc
          6845 => x"84", -- $01abd
          6846 => x"83", -- $01abe
          6847 => x"82", -- $01abf
          6848 => x"82", -- $01ac0
          6849 => x"81", -- $01ac1
          6850 => x"81", -- $01ac2
          6851 => x"81", -- $01ac3
          6852 => x"80", -- $01ac4
          6853 => x"80", -- $01ac5
          6854 => x"80", -- $01ac6
          6855 => x"80", -- $01ac7
          6856 => x"80", -- $01ac8
          6857 => x"80", -- $01ac9
          6858 => x"81", -- $01aca
          6859 => x"82", -- $01acb
          6860 => x"83", -- $01acc
          6861 => x"83", -- $01acd
          6862 => x"84", -- $01ace
          6863 => x"84", -- $01acf
          6864 => x"83", -- $01ad0
          6865 => x"82", -- $01ad1
          6866 => x"81", -- $01ad2
          6867 => x"80", -- $01ad3
          6868 => x"80", -- $01ad4
          6869 => x"80", -- $01ad5
          6870 => x"7f", -- $01ad6
          6871 => x"7f", -- $01ad7
          6872 => x"80", -- $01ad8
          6873 => x"80", -- $01ad9
          6874 => x"82", -- $01ada
          6875 => x"84", -- $01adb
          6876 => x"85", -- $01adc
          6877 => x"86", -- $01add
          6878 => x"87", -- $01ade
          6879 => x"87", -- $01adf
          6880 => x"85", -- $01ae0
          6881 => x"84", -- $01ae1
          6882 => x"83", -- $01ae2
          6883 => x"80", -- $01ae3
          6884 => x"80", -- $01ae4
          6885 => x"7f", -- $01ae5
          6886 => x"7f", -- $01ae6
          6887 => x"7f", -- $01ae7
          6888 => x"80", -- $01ae8
          6889 => x"83", -- $01ae9
          6890 => x"85", -- $01aea
          6891 => x"87", -- $01aeb
          6892 => x"88", -- $01aec
          6893 => x"88", -- $01aed
          6894 => x"88", -- $01aee
          6895 => x"88", -- $01aef
          6896 => x"88", -- $01af0
          6897 => x"88", -- $01af1
          6898 => x"88", -- $01af2
          6899 => x"87", -- $01af3
          6900 => x"86", -- $01af4
          6901 => x"84", -- $01af5
          6902 => x"83", -- $01af6
          6903 => x"81", -- $01af7
          6904 => x"80", -- $01af8
          6905 => x"80", -- $01af9
          6906 => x"80", -- $01afa
          6907 => x"80", -- $01afb
          6908 => x"81", -- $01afc
          6909 => x"81", -- $01afd
          6910 => x"80", -- $01afe
          6911 => x"80", -- $01aff
          6912 => x"7e", -- $01b00
          6913 => x"7b", -- $01b01
          6914 => x"79", -- $01b02
          6915 => x"78", -- $01b03
          6916 => x"77", -- $01b04
          6917 => x"78", -- $01b05
          6918 => x"7a", -- $01b06
          6919 => x"7d", -- $01b07
          6920 => x"80", -- $01b08
          6921 => x"82", -- $01b09
          6922 => x"83", -- $01b0a
          6923 => x"84", -- $01b0b
          6924 => x"85", -- $01b0c
          6925 => x"84", -- $01b0d
          6926 => x"84", -- $01b0e
          6927 => x"83", -- $01b0f
          6928 => x"83", -- $01b10
          6929 => x"82", -- $01b11
          6930 => x"82", -- $01b12
          6931 => x"82", -- $01b13
          6932 => x"81", -- $01b14
          6933 => x"80", -- $01b15
          6934 => x"80", -- $01b16
          6935 => x"7f", -- $01b17
          6936 => x"7e", -- $01b18
          6937 => x"7e", -- $01b19
          6938 => x"7e", -- $01b1a
          6939 => x"7e", -- $01b1b
          6940 => x"7f", -- $01b1c
          6941 => x"80", -- $01b1d
          6942 => x"80", -- $01b1e
          6943 => x"81", -- $01b1f
          6944 => x"82", -- $01b20
          6945 => x"82", -- $01b21
          6946 => x"83", -- $01b22
          6947 => x"82", -- $01b23
          6948 => x"82", -- $01b24
          6949 => x"81", -- $01b25
          6950 => x"81", -- $01b26
          6951 => x"81", -- $01b27
          6952 => x"81", -- $01b28
          6953 => x"81", -- $01b29
          6954 => x"81", -- $01b2a
          6955 => x"82", -- $01b2b
          6956 => x"82", -- $01b2c
          6957 => x"82", -- $01b2d
          6958 => x"82", -- $01b2e
          6959 => x"82", -- $01b2f
          6960 => x"82", -- $01b30
          6961 => x"82", -- $01b31
          6962 => x"82", -- $01b32
          6963 => x"82", -- $01b33
          6964 => x"82", -- $01b34
          6965 => x"82", -- $01b35
          6966 => x"82", -- $01b36
          6967 => x"83", -- $01b37
          6968 => x"84", -- $01b38
          6969 => x"85", -- $01b39
          6970 => x"86", -- $01b3a
          6971 => x"87", -- $01b3b
          6972 => x"87", -- $01b3c
          6973 => x"87", -- $01b3d
          6974 => x"85", -- $01b3e
          6975 => x"84", -- $01b3f
          6976 => x"82", -- $01b40
          6977 => x"80", -- $01b41
          6978 => x"80", -- $01b42
          6979 => x"80", -- $01b43
          6980 => x"80", -- $01b44
          6981 => x"81", -- $01b45
          6982 => x"82", -- $01b46
          6983 => x"82", -- $01b47
          6984 => x"82", -- $01b48
          6985 => x"80", -- $01b49
          6986 => x"7e", -- $01b4a
          6987 => x"7b", -- $01b4b
          6988 => x"78", -- $01b4c
          6989 => x"76", -- $01b4d
          6990 => x"75", -- $01b4e
          6991 => x"75", -- $01b4f
          6992 => x"77", -- $01b50
          6993 => x"79", -- $01b51
          6994 => x"7b", -- $01b52
          6995 => x"7e", -- $01b53
          6996 => x"80", -- $01b54
          6997 => x"81", -- $01b55
          6998 => x"82", -- $01b56
          6999 => x"82", -- $01b57
          7000 => x"81", -- $01b58
          7001 => x"81", -- $01b59
          7002 => x"80", -- $01b5a
          7003 => x"80", -- $01b5b
          7004 => x"80", -- $01b5c
          7005 => x"80", -- $01b5d
          7006 => x"80", -- $01b5e
          7007 => x"80", -- $01b5f
          7008 => x"80", -- $01b60
          7009 => x"80", -- $01b61
          7010 => x"80", -- $01b62
          7011 => x"7f", -- $01b63
          7012 => x"7f", -- $01b64
          7013 => x"7f", -- $01b65
          7014 => x"7f", -- $01b66
          7015 => x"7f", -- $01b67
          7016 => x"80", -- $01b68
          7017 => x"80", -- $01b69
          7018 => x"80", -- $01b6a
          7019 => x"80", -- $01b6b
          7020 => x"80", -- $01b6c
          7021 => x"80", -- $01b6d
          7022 => x"80", -- $01b6e
          7023 => x"80", -- $01b6f
          7024 => x"80", -- $01b70
          7025 => x"80", -- $01b71
          7026 => x"80", -- $01b72
          7027 => x"80", -- $01b73
          7028 => x"80", -- $01b74
          7029 => x"81", -- $01b75
          7030 => x"81", -- $01b76
          7031 => x"82", -- $01b77
          7032 => x"83", -- $01b78
          7033 => x"83", -- $01b79
          7034 => x"83", -- $01b7a
          7035 => x"83", -- $01b7b
          7036 => x"82", -- $01b7c
          7037 => x"82", -- $01b7d
          7038 => x"81", -- $01b7e
          7039 => x"81", -- $01b7f
          7040 => x"80", -- $01b80
          7041 => x"80", -- $01b81
          7042 => x"81", -- $01b82
          7043 => x"81", -- $01b83
          7044 => x"82", -- $01b84
          7045 => x"83", -- $01b85
          7046 => x"84", -- $01b86
          7047 => x"85", -- $01b87
          7048 => x"86", -- $01b88
          7049 => x"86", -- $01b89
          7050 => x"86", -- $01b8a
          7051 => x"85", -- $01b8b
          7052 => x"83", -- $01b8c
          7053 => x"81", -- $01b8d
          7054 => x"80", -- $01b8e
          7055 => x"80", -- $01b8f
          7056 => x"80", -- $01b90
          7057 => x"80", -- $01b91
          7058 => x"80", -- $01b92
          7059 => x"80", -- $01b93
          7060 => x"80", -- $01b94
          7061 => x"7f", -- $01b95
          7062 => x"7d", -- $01b96
          7063 => x"7c", -- $01b97
          7064 => x"7a", -- $01b98
          7065 => x"79", -- $01b99
          7066 => x"78", -- $01b9a
          7067 => x"77", -- $01b9b
          7068 => x"78", -- $01b9c
          7069 => x"7a", -- $01b9d
          7070 => x"7b", -- $01b9e
          7071 => x"7c", -- $01b9f
          7072 => x"7e", -- $01ba0
          7073 => x"7f", -- $01ba1
          7074 => x"7f", -- $01ba2
          7075 => x"80", -- $01ba3
          7076 => x"80", -- $01ba4
          7077 => x"80", -- $01ba5
          7078 => x"80", -- $01ba6
          7079 => x"80", -- $01ba7
          7080 => x"80", -- $01ba8
          7081 => x"80", -- $01ba9
          7082 => x"80", -- $01baa
          7083 => x"80", -- $01bab
          7084 => x"80", -- $01bac
          7085 => x"80", -- $01bad
          7086 => x"80", -- $01bae
          7087 => x"80", -- $01baf
          7088 => x"80", -- $01bb0
          7089 => x"80", -- $01bb1
          7090 => x"7f", -- $01bb2
          7091 => x"7f", -- $01bb3
          7092 => x"7f", -- $01bb4
          7093 => x"7f", -- $01bb5
          7094 => x"80", -- $01bb6
          7095 => x"80", -- $01bb7
          7096 => x"80", -- $01bb8
          7097 => x"80", -- $01bb9
          7098 => x"80", -- $01bba
          7099 => x"80", -- $01bbb
          7100 => x"80", -- $01bbc
          7101 => x"80", -- $01bbd
          7102 => x"80", -- $01bbe
          7103 => x"80", -- $01bbf
          7104 => x"80", -- $01bc0
          7105 => x"80", -- $01bc1
          7106 => x"80", -- $01bc2
          7107 => x"80", -- $01bc3
          7108 => x"81", -- $01bc4
          7109 => x"81", -- $01bc5
          7110 => x"81", -- $01bc6
          7111 => x"81", -- $01bc7
          7112 => x"80", -- $01bc8
          7113 => x"80", -- $01bc9
          7114 => x"80", -- $01bca
          7115 => x"80", -- $01bcb
          7116 => x"7f", -- $01bcc
          7117 => x"7e", -- $01bcd
          7118 => x"7f", -- $01bce
          7119 => x"7f", -- $01bcf
          7120 => x"7f", -- $01bd0
          7121 => x"80", -- $01bd1
          7122 => x"80", -- $01bd2
          7123 => x"81", -- $01bd3
          7124 => x"82", -- $01bd4
          7125 => x"84", -- $01bd5
          7126 => x"84", -- $01bd6
          7127 => x"84", -- $01bd7
          7128 => x"84", -- $01bd8
          7129 => x"83", -- $01bd9
          7130 => x"82", -- $01bda
          7131 => x"81", -- $01bdb
          7132 => x"81", -- $01bdc
          7133 => x"81", -- $01bdd
          7134 => x"80", -- $01bde
          7135 => x"80", -- $01bdf
          7136 => x"80", -- $01be0
          7137 => x"80", -- $01be1
          7138 => x"7f", -- $01be2
          7139 => x"7e", -- $01be3
          7140 => x"7c", -- $01be4
          7141 => x"7b", -- $01be5
          7142 => x"79", -- $01be6
          7143 => x"78", -- $01be7
          7144 => x"77", -- $01be8
          7145 => x"77", -- $01be9
          7146 => x"76", -- $01bea
          7147 => x"77", -- $01beb
          7148 => x"78", -- $01bec
          7149 => x"78", -- $01bed
          7150 => x"79", -- $01bee
          7151 => x"7a", -- $01bef
          7152 => x"7b", -- $01bf0
          7153 => x"7c", -- $01bf1
          7154 => x"7d", -- $01bf2
          7155 => x"7f", -- $01bf3
          7156 => x"80", -- $01bf4
          7157 => x"80", -- $01bf5
          7158 => x"81", -- $01bf6
          7159 => x"82", -- $01bf7
          7160 => x"82", -- $01bf8
          7161 => x"82", -- $01bf9
          7162 => x"82", -- $01bfa
          7163 => x"81", -- $01bfb
          7164 => x"80", -- $01bfc
          7165 => x"80", -- $01bfd
          7166 => x"7f", -- $01bfe
          7167 => x"7d", -- $01bff
          7168 => x"7d", -- $01c00
          7169 => x"7c", -- $01c01
          7170 => x"7b", -- $01c02
          7171 => x"7b", -- $01c03
          7172 => x"7b", -- $01c04
          7173 => x"7c", -- $01c05
          7174 => x"7d", -- $01c06
          7175 => x"7e", -- $01c07
          7176 => x"7e", -- $01c08
          7177 => x"7f", -- $01c09
          7178 => x"7f", -- $01c0a
          7179 => x"7f", -- $01c0b
          7180 => x"7f", -- $01c0c
          7181 => x"7f", -- $01c0d
          7182 => x"7e", -- $01c0e
          7183 => x"7e", -- $01c0f
          7184 => x"7e", -- $01c10
          7185 => x"7e", -- $01c11
          7186 => x"7f", -- $01c12
          7187 => x"7f", -- $01c13
          7188 => x"7f", -- $01c14
          7189 => x"7f", -- $01c15
          7190 => x"80", -- $01c16
          7191 => x"80", -- $01c17
          7192 => x"80", -- $01c18
          7193 => x"80", -- $01c19
          7194 => x"80", -- $01c1a
          7195 => x"80", -- $01c1b
          7196 => x"80", -- $01c1c
          7197 => x"80", -- $01c1d
          7198 => x"80", -- $01c1e
          7199 => x"80", -- $01c1f
          7200 => x"80", -- $01c20
          7201 => x"80", -- $01c21
          7202 => x"80", -- $01c22
          7203 => x"80", -- $01c23
          7204 => x"81", -- $01c24
          7205 => x"81", -- $01c25
          7206 => x"81", -- $01c26
          7207 => x"81", -- $01c27
          7208 => x"81", -- $01c28
          7209 => x"81", -- $01c29
          7210 => x"82", -- $01c2a
          7211 => x"81", -- $01c2b
          7212 => x"81", -- $01c2c
          7213 => x"81", -- $01c2d
          7214 => x"80", -- $01c2e
          7215 => x"80", -- $01c2f
          7216 => x"7f", -- $01c30
          7217 => x"7d", -- $01c31
          7218 => x"7c", -- $01c32
          7219 => x"7b", -- $01c33
          7220 => x"7a", -- $01c34
          7221 => x"79", -- $01c35
          7222 => x"79", -- $01c36
          7223 => x"79", -- $01c37
          7224 => x"79", -- $01c38
          7225 => x"79", -- $01c39
          7226 => x"79", -- $01c3a
          7227 => x"79", -- $01c3b
          7228 => x"79", -- $01c3c
          7229 => x"7a", -- $01c3d
          7230 => x"7a", -- $01c3e
          7231 => x"7b", -- $01c3f
          7232 => x"7c", -- $01c40
          7233 => x"7c", -- $01c41
          7234 => x"7d", -- $01c42
          7235 => x"7e", -- $01c43
          7236 => x"7e", -- $01c44
          7237 => x"7f", -- $01c45
          7238 => x"80", -- $01c46
          7239 => x"80", -- $01c47
          7240 => x"80", -- $01c48
          7241 => x"81", -- $01c49
          7242 => x"81", -- $01c4a
          7243 => x"81", -- $01c4b
          7244 => x"81", -- $01c4c
          7245 => x"81", -- $01c4d
          7246 => x"80", -- $01c4e
          7247 => x"80", -- $01c4f
          7248 => x"80", -- $01c50
          7249 => x"7f", -- $01c51
          7250 => x"7e", -- $01c52
          7251 => x"7e", -- $01c53
          7252 => x"7e", -- $01c54
          7253 => x"7d", -- $01c55
          7254 => x"7d", -- $01c56
          7255 => x"7d", -- $01c57
          7256 => x"7d", -- $01c58
          7257 => x"7d", -- $01c59
          7258 => x"7e", -- $01c5a
          7259 => x"7e", -- $01c5b
          7260 => x"7f", -- $01c5c
          7261 => x"7f", -- $01c5d
          7262 => x"7f", -- $01c5e
          7263 => x"80", -- $01c5f
          7264 => x"80", -- $01c60
          7265 => x"80", -- $01c61
          7266 => x"80", -- $01c62
          7267 => x"80", -- $01c63
          7268 => x"7f", -- $01c64
          7269 => x"7f", -- $01c65
          7270 => x"7f", -- $01c66
          7271 => x"7f", -- $01c67
          7272 => x"7f", -- $01c68
          7273 => x"80", -- $01c69
          7274 => x"80", -- $01c6a
          7275 => x"80", -- $01c6b
          7276 => x"80", -- $01c6c
          7277 => x"80", -- $01c6d
          7278 => x"81", -- $01c6e
          7279 => x"82", -- $01c6f
          7280 => x"82", -- $01c70
          7281 => x"83", -- $01c71
          7282 => x"83", -- $01c72
          7283 => x"83", -- $01c73
          7284 => x"83", -- $01c74
          7285 => x"83", -- $01c75
          7286 => x"82", -- $01c76
          7287 => x"82", -- $01c77
          7288 => x"81", -- $01c78
          7289 => x"80", -- $01c79
          7290 => x"80", -- $01c7a
          7291 => x"80", -- $01c7b
          7292 => x"80", -- $01c7c
          7293 => x"80", -- $01c7d
          7294 => x"80", -- $01c7e
          7295 => x"80", -- $01c7f
          7296 => x"80", -- $01c80
          7297 => x"7f", -- $01c81
          7298 => x"7e", -- $01c82
          7299 => x"7d", -- $01c83
          7300 => x"7d", -- $01c84
          7301 => x"7d", -- $01c85
          7302 => x"7c", -- $01c86
          7303 => x"7b", -- $01c87
          7304 => x"7b", -- $01c88
          7305 => x"7a", -- $01c89
          7306 => x"7a", -- $01c8a
          7307 => x"7a", -- $01c8b
          7308 => x"7a", -- $01c8c
          7309 => x"7a", -- $01c8d
          7310 => x"7b", -- $01c8e
          7311 => x"7b", -- $01c8f
          7312 => x"7c", -- $01c90
          7313 => x"7d", -- $01c91
          7314 => x"7e", -- $01c92
          7315 => x"7e", -- $01c93
          7316 => x"7f", -- $01c94
          7317 => x"7f", -- $01c95
          7318 => x"7f", -- $01c96
          7319 => x"7f", -- $01c97
          7320 => x"7f", -- $01c98
          7321 => x"7f", -- $01c99
          7322 => x"7f", -- $01c9a
          7323 => x"7f", -- $01c9b
          7324 => x"7f", -- $01c9c
          7325 => x"7f", -- $01c9d
          7326 => x"7f", -- $01c9e
          7327 => x"7f", -- $01c9f
          7328 => x"7f", -- $01ca0
          7329 => x"7f", -- $01ca1
          7330 => x"80", -- $01ca2
          7331 => x"80", -- $01ca3
          7332 => x"80", -- $01ca4
          7333 => x"80", -- $01ca5
          7334 => x"80", -- $01ca6
          7335 => x"80", -- $01ca7
          7336 => x"80", -- $01ca8
          7337 => x"80", -- $01ca9
          7338 => x"80", -- $01caa
          7339 => x"80", -- $01cab
          7340 => x"80", -- $01cac
          7341 => x"80", -- $01cad
          7342 => x"80", -- $01cae
          7343 => x"80", -- $01caf
          7344 => x"80", -- $01cb0
          7345 => x"80", -- $01cb1
          7346 => x"80", -- $01cb2
          7347 => x"80", -- $01cb3
          7348 => x"80", -- $01cb4
          7349 => x"80", -- $01cb5
          7350 => x"80", -- $01cb6
          7351 => x"80", -- $01cb7
          7352 => x"80", -- $01cb8
          7353 => x"80", -- $01cb9
          7354 => x"80", -- $01cba
          7355 => x"81", -- $01cbb
          7356 => x"81", -- $01cbc
          7357 => x"82", -- $01cbd
          7358 => x"82", -- $01cbe
          7359 => x"83", -- $01cbf
          7360 => x"83", -- $01cc0
          7361 => x"83", -- $01cc1
          7362 => x"83", -- $01cc2
          7363 => x"84", -- $01cc3
          7364 => x"84", -- $01cc4
          7365 => x"84", -- $01cc5
          7366 => x"84", -- $01cc6
          7367 => x"83", -- $01cc7
          7368 => x"83", -- $01cc8
          7369 => x"82", -- $01cc9
          7370 => x"80", -- $01cca
          7371 => x"80", -- $01ccb
          7372 => x"7f", -- $01ccc
          7373 => x"7d", -- $01ccd
          7374 => x"7c", -- $01cce
          7375 => x"7b", -- $01ccf
          7376 => x"7a", -- $01cd0
          7377 => x"7a", -- $01cd1
          7378 => x"79", -- $01cd2
          7379 => x"78", -- $01cd3
          7380 => x"78", -- $01cd4
          7381 => x"77", -- $01cd5
          7382 => x"78", -- $01cd6
          7383 => x"78", -- $01cd7
          7384 => x"78", -- $01cd8
          7385 => x"78", -- $01cd9
          7386 => x"7a", -- $01cda
          7387 => x"7b", -- $01cdb
          7388 => x"7c", -- $01cdc
          7389 => x"7d", -- $01cdd
          7390 => x"7e", -- $01cde
          7391 => x"7f", -- $01cdf
          7392 => x"80", -- $01ce0
          7393 => x"80", -- $01ce1
          7394 => x"81", -- $01ce2
          7395 => x"81", -- $01ce3
          7396 => x"81", -- $01ce4
          7397 => x"82", -- $01ce5
          7398 => x"82", -- $01ce6
          7399 => x"82", -- $01ce7
          7400 => x"82", -- $01ce8
          7401 => x"81", -- $01ce9
          7402 => x"81", -- $01cea
          7403 => x"80", -- $01ceb
          7404 => x"80", -- $01cec
          7405 => x"80", -- $01ced
          7406 => x"80", -- $01cee
          7407 => x"80", -- $01cef
          7408 => x"80", -- $01cf0
          7409 => x"80", -- $01cf1
          7410 => x"80", -- $01cf2
          7411 => x"80", -- $01cf3
          7412 => x"80", -- $01cf4
          7413 => x"80", -- $01cf5
          7414 => x"80", -- $01cf6
          7415 => x"80", -- $01cf7
          7416 => x"80", -- $01cf8
          7417 => x"80", -- $01cf9
          7418 => x"80", -- $01cfa
          7419 => x"80", -- $01cfb
          7420 => x"80", -- $01cfc
          7421 => x"80", -- $01cfd
          7422 => x"80", -- $01cfe
          7423 => x"80", -- $01cff
          7424 => x"80", -- $01d00
          7425 => x"80", -- $01d01
          7426 => x"80", -- $01d02
          7427 => x"80", -- $01d03
          7428 => x"80", -- $01d04
          7429 => x"81", -- $01d05
          7430 => x"81", -- $01d06
          7431 => x"81", -- $01d07
          7432 => x"82", -- $01d08
          7433 => x"82", -- $01d09
          7434 => x"83", -- $01d0a
          7435 => x"83", -- $01d0b
          7436 => x"83", -- $01d0c
          7437 => x"83", -- $01d0d
          7438 => x"83", -- $01d0e
          7439 => x"84", -- $01d0f
          7440 => x"84", -- $01d10
          7441 => x"83", -- $01d11
          7442 => x"83", -- $01d12
          7443 => x"83", -- $01d13
          7444 => x"83", -- $01d14
          7445 => x"83", -- $01d15
          7446 => x"82", -- $01d16
          7447 => x"82", -- $01d17
          7448 => x"81", -- $01d18
          7449 => x"81", -- $01d19
          7450 => x"80", -- $01d1a
          7451 => x"80", -- $01d1b
          7452 => x"80", -- $01d1c
          7453 => x"7f", -- $01d1d
          7454 => x"7e", -- $01d1e
          7455 => x"7d", -- $01d1f
          7456 => x"7c", -- $01d20
          7457 => x"7b", -- $01d21
          7458 => x"7a", -- $01d22
          7459 => x"7a", -- $01d23
          7460 => x"7a", -- $01d24
          7461 => x"79", -- $01d25
          7462 => x"79", -- $01d26
          7463 => x"7a", -- $01d27
          7464 => x"7a", -- $01d28
          7465 => x"7b", -- $01d29
          7466 => x"7b", -- $01d2a
          7467 => x"7c", -- $01d2b
          7468 => x"7e", -- $01d2c
          7469 => x"7e", -- $01d2d
          7470 => x"7f", -- $01d2e
          7471 => x"80", -- $01d2f
          7472 => x"80", -- $01d30
          7473 => x"80", -- $01d31
          7474 => x"81", -- $01d32
          7475 => x"81", -- $01d33
          7476 => x"82", -- $01d34
          7477 => x"82", -- $01d35
          7478 => x"82", -- $01d36
          7479 => x"82", -- $01d37
          7480 => x"82", -- $01d38
          7481 => x"82", -- $01d39
          7482 => x"82", -- $01d3a
          7483 => x"82", -- $01d3b
          7484 => x"82", -- $01d3c
          7485 => x"82", -- $01d3d
          7486 => x"82", -- $01d3e
          7487 => x"82", -- $01d3f
          7488 => x"82", -- $01d40
          7489 => x"82", -- $01d41
          7490 => x"82", -- $01d42
          7491 => x"82", -- $01d43
          7492 => x"81", -- $01d44
          7493 => x"81", -- $01d45
          7494 => x"81", -- $01d46
          7495 => x"80", -- $01d47
          7496 => x"80", -- $01d48
          7497 => x"80", -- $01d49
          7498 => x"80", -- $01d4a
          7499 => x"80", -- $01d4b
          7500 => x"80", -- $01d4c
          7501 => x"80", -- $01d4d
          7502 => x"80", -- $01d4e
          7503 => x"81", -- $01d4f
          7504 => x"81", -- $01d50
          7505 => x"81", -- $01d51
          7506 => x"82", -- $01d52
          7507 => x"82", -- $01d53
          7508 => x"83", -- $01d54
          7509 => x"83", -- $01d55
          7510 => x"83", -- $01d56
          7511 => x"84", -- $01d57
          7512 => x"84", -- $01d58
          7513 => x"84", -- $01d59
          7514 => x"84", -- $01d5a
          7515 => x"83", -- $01d5b
          7516 => x"83", -- $01d5c
          7517 => x"83", -- $01d5d
          7518 => x"84", -- $01d5e
          7519 => x"84", -- $01d5f
          7520 => x"84", -- $01d60
          7521 => x"84", -- $01d61
          7522 => x"84", -- $01d62
          7523 => x"84", -- $01d63
          7524 => x"83", -- $01d64
          7525 => x"83", -- $01d65
          7526 => x"82", -- $01d66
          7527 => x"82", -- $01d67
          7528 => x"81", -- $01d68
          7529 => x"81", -- $01d69
          7530 => x"80", -- $01d6a
          7531 => x"80", -- $01d6b
          7532 => x"7f", -- $01d6c
          7533 => x"7e", -- $01d6d
          7534 => x"7e", -- $01d6e
          7535 => x"7d", -- $01d6f
          7536 => x"7c", -- $01d70
          7537 => x"7c", -- $01d71
          7538 => x"7c", -- $01d72
          7539 => x"7c", -- $01d73
          7540 => x"7c", -- $01d74
          7541 => x"7c", -- $01d75
          7542 => x"7d", -- $01d76
          7543 => x"7d", -- $01d77
          7544 => x"7e", -- $01d78
          7545 => x"7f", -- $01d79
          7546 => x"7f", -- $01d7a
          7547 => x"80", -- $01d7b
          7548 => x"80", -- $01d7c
          7549 => x"80", -- $01d7d
          7550 => x"80", -- $01d7e
          7551 => x"81", -- $01d7f
          7552 => x"81", -- $01d80
          7553 => x"81", -- $01d81
          7554 => x"82", -- $01d82
          7555 => x"82", -- $01d83
          7556 => x"82", -- $01d84
          7557 => x"82", -- $01d85
          7558 => x"83", -- $01d86
          7559 => x"83", -- $01d87
          7560 => x"83", -- $01d88
          7561 => x"83", -- $01d89
          7562 => x"83", -- $01d8a
          7563 => x"82", -- $01d8b
          7564 => x"82", -- $01d8c
          7565 => x"82", -- $01d8d
          7566 => x"81", -- $01d8e
          7567 => x"81", -- $01d8f
          7568 => x"81", -- $01d90
          7569 => x"81", -- $01d91
          7570 => x"81", -- $01d92
          7571 => x"81", -- $01d93
          7572 => x"81", -- $01d94
          7573 => x"81", -- $01d95
          7574 => x"81", -- $01d96
          7575 => x"81", -- $01d97
          7576 => x"81", -- $01d98
          7577 => x"80", -- $01d99
          7578 => x"80", -- $01d9a
          7579 => x"80", -- $01d9b
          7580 => x"80", -- $01d9c
          7581 => x"80", -- $01d9d
          7582 => x"80", -- $01d9e
          7583 => x"80", -- $01d9f
          7584 => x"80", -- $01da0
          7585 => x"80", -- $01da1
          7586 => x"80", -- $01da2
          7587 => x"80", -- $01da3
          7588 => x"80", -- $01da4
          7589 => x"80", -- $01da5
          7590 => x"81", -- $01da6
          7591 => x"81", -- $01da7
          7592 => x"81", -- $01da8
          7593 => x"82", -- $01da9
          7594 => x"83", -- $01daa
          7595 => x"83", -- $01dab
          7596 => x"84", -- $01dac
          7597 => x"84", -- $01dad
          7598 => x"84", -- $01dae
          7599 => x"84", -- $01daf
          7600 => x"84", -- $01db0
          7601 => x"84", -- $01db1
          7602 => x"84", -- $01db2
          7603 => x"84", -- $01db3
          7604 => x"83", -- $01db4
          7605 => x"82", -- $01db5
          7606 => x"82", -- $01db6
          7607 => x"81", -- $01db7
          7608 => x"80", -- $01db8
          7609 => x"80", -- $01db9
          7610 => x"7f", -- $01dba
          7611 => x"7e", -- $01dbb
          7612 => x"7d", -- $01dbc
          7613 => x"7c", -- $01dbd
          7614 => x"7b", -- $01dbe
          7615 => x"7b", -- $01dbf
          7616 => x"7a", -- $01dc0
          7617 => x"7a", -- $01dc1
          7618 => x"7a", -- $01dc2
          7619 => x"7a", -- $01dc3
          7620 => x"7a", -- $01dc4
          7621 => x"7b", -- $01dc5
          7622 => x"7b", -- $01dc6
          7623 => x"7c", -- $01dc7
          7624 => x"7c", -- $01dc8
          7625 => x"7d", -- $01dc9
          7626 => x"7e", -- $01dca
          7627 => x"7f", -- $01dcb
          7628 => x"80", -- $01dcc
          7629 => x"80", -- $01dcd
          7630 => x"80", -- $01dce
          7631 => x"81", -- $01dcf
          7632 => x"82", -- $01dd0
          7633 => x"82", -- $01dd1
          7634 => x"83", -- $01dd2
          7635 => x"83", -- $01dd3
          7636 => x"83", -- $01dd4
          7637 => x"83", -- $01dd5
          7638 => x"83", -- $01dd6
          7639 => x"83", -- $01dd7
          7640 => x"83", -- $01dd8
          7641 => x"82", -- $01dd9
          7642 => x"82", -- $01dda
          7643 => x"82", -- $01ddb
          7644 => x"82", -- $01ddc
          7645 => x"81", -- $01ddd
          7646 => x"82", -- $01dde
          7647 => x"81", -- $01ddf
          7648 => x"81", -- $01de0
          7649 => x"81", -- $01de1
          7650 => x"81", -- $01de2
          7651 => x"81", -- $01de3
          7652 => x"81", -- $01de4
          7653 => x"81", -- $01de5
          7654 => x"80", -- $01de6
          7655 => x"80", -- $01de7
          7656 => x"80", -- $01de8
          7657 => x"80", -- $01de9
          7658 => x"80", -- $01dea
          7659 => x"80", -- $01deb
          7660 => x"80", -- $01dec
          7661 => x"80", -- $01ded
          7662 => x"80", -- $01dee
          7663 => x"80", -- $01def
          7664 => x"80", -- $01df0
          7665 => x"80", -- $01df1
          7666 => x"80", -- $01df2
          7667 => x"81", -- $01df3
          7668 => x"81", -- $01df4
          7669 => x"82", -- $01df5
          7670 => x"82", -- $01df6
          7671 => x"83", -- $01df7
          7672 => x"83", -- $01df8
          7673 => x"83", -- $01df9
          7674 => x"84", -- $01dfa
          7675 => x"84", -- $01dfb
          7676 => x"84", -- $01dfc
          7677 => x"85", -- $01dfd
          7678 => x"85", -- $01dfe
          7679 => x"85", -- $01dff
          7680 => x"85", -- $01e00
          7681 => x"84", -- $01e01
          7682 => x"84", -- $01e02
          7683 => x"83", -- $01e03
          7684 => x"83", -- $01e04
          7685 => x"82", -- $01e05
          7686 => x"81", -- $01e06
          7687 => x"80", -- $01e07
          7688 => x"80", -- $01e08
          7689 => x"7f", -- $01e09
          7690 => x"7e", -- $01e0a
          7691 => x"7d", -- $01e0b
          7692 => x"7d", -- $01e0c
          7693 => x"7c", -- $01e0d
          7694 => x"7b", -- $01e0e
          7695 => x"7b", -- $01e0f
          7696 => x"7b", -- $01e10
          7697 => x"7b", -- $01e11
          7698 => x"7b", -- $01e12
          7699 => x"7c", -- $01e13
          7700 => x"7c", -- $01e14
          7701 => x"7d", -- $01e15
          7702 => x"7d", -- $01e16
          7703 => x"7e", -- $01e17
          7704 => x"7f", -- $01e18
          7705 => x"80", -- $01e19
          7706 => x"80", -- $01e1a
          7707 => x"80", -- $01e1b
          7708 => x"81", -- $01e1c
          7709 => x"82", -- $01e1d
          7710 => x"83", -- $01e1e
          7711 => x"83", -- $01e1f
          7712 => x"84", -- $01e20
          7713 => x"84", -- $01e21
          7714 => x"84", -- $01e22
          7715 => x"85", -- $01e23
          7716 => x"85", -- $01e24
          7717 => x"85", -- $01e25
          7718 => x"85", -- $01e26
          7719 => x"84", -- $01e27
          7720 => x"84", -- $01e28
          7721 => x"84", -- $01e29
          7722 => x"84", -- $01e2a
          7723 => x"83", -- $01e2b
          7724 => x"83", -- $01e2c
          7725 => x"83", -- $01e2d
          7726 => x"82", -- $01e2e
          7727 => x"82", -- $01e2f
          7728 => x"82", -- $01e30
          7729 => x"81", -- $01e31
          7730 => x"81", -- $01e32
          7731 => x"80", -- $01e33
          7732 => x"80", -- $01e34
          7733 => x"80", -- $01e35
          7734 => x"80", -- $01e36
          7735 => x"80", -- $01e37
          7736 => x"80", -- $01e38
          7737 => x"80", -- $01e39
          7738 => x"80", -- $01e3a
          7739 => x"80", -- $01e3b
          7740 => x"80", -- $01e3c
          7741 => x"80", -- $01e3d
          7742 => x"81", -- $01e3e
          7743 => x"81", -- $01e3f
          7744 => x"82", -- $01e40
          7745 => x"82", -- $01e41
          7746 => x"82", -- $01e42
          7747 => x"83", -- $01e43
          7748 => x"83", -- $01e44
          7749 => x"83", -- $01e45
          7750 => x"84", -- $01e46
          7751 => x"84", -- $01e47
          7752 => x"83", -- $01e48
          7753 => x"84", -- $01e49
          7754 => x"84", -- $01e4a
          7755 => x"84", -- $01e4b
          7756 => x"84", -- $01e4c
          7757 => x"84", -- $01e4d
          7758 => x"83", -- $01e4e
          7759 => x"82", -- $01e4f
          7760 => x"82", -- $01e50
          7761 => x"81", -- $01e51
          7762 => x"80", -- $01e52
          7763 => x"80", -- $01e53
          7764 => x"7f", -- $01e54
          7765 => x"7e", -- $01e55
          7766 => x"7e", -- $01e56
          7767 => x"79", -- $01e57
          7768 => x"77", -- $01e58
          7769 => x"77", -- $01e59
          7770 => x"79", -- $01e5a
          7771 => x"7a", -- $01e5b
          7772 => x"7a", -- $01e5c
          7773 => x"7a", -- $01e5d
          7774 => x"7a", -- $01e5e
          7775 => x"7a", -- $01e5f
          7776 => x"7a", -- $01e60
          7777 => x"7a", -- $01e61
          7778 => x"7b", -- $01e62
          7779 => x"7b", -- $01e63
          7780 => x"7c", -- $01e64
          7781 => x"7e", -- $01e65
          7782 => x"7f", -- $01e66
          7783 => x"80", -- $01e67
          7784 => x"82", -- $01e68
          7785 => x"83", -- $01e69
          7786 => x"85", -- $01e6a
          7787 => x"86", -- $01e6b
          7788 => x"86", -- $01e6c
          7789 => x"85", -- $01e6d
          7790 => x"85", -- $01e6e
          7791 => x"85", -- $01e6f
          7792 => x"84", -- $01e70
          7793 => x"84", -- $01e71
          7794 => x"83", -- $01e72
          7795 => x"82", -- $01e73
          7796 => x"80", -- $01e74
          7797 => x"80", -- $01e75
          7798 => x"80", -- $01e76
          7799 => x"7f", -- $01e77
          7800 => x"7f", -- $01e78
          7801 => x"7f", -- $01e79
          7802 => x"7f", -- $01e7a
          7803 => x"7f", -- $01e7b
          7804 => x"7f", -- $01e7c
          7805 => x"7f", -- $01e7d
          7806 => x"7f", -- $01e7e
          7807 => x"7f", -- $01e7f
          7808 => x"80", -- $01e80
          7809 => x"80", -- $01e81
          7810 => x"80", -- $01e82
          7811 => x"81", -- $01e83
          7812 => x"81", -- $01e84
          7813 => x"81", -- $01e85
          7814 => x"80", -- $01e86
          7815 => x"80", -- $01e87
          7816 => x"80", -- $01e88
          7817 => x"80", -- $01e89
          7818 => x"80", -- $01e8a
          7819 => x"81", -- $01e8b
          7820 => x"82", -- $01e8c
          7821 => x"84", -- $01e8d
          7822 => x"84", -- $01e8e
          7823 => x"84", -- $01e8f
          7824 => x"83", -- $01e90
          7825 => x"83", -- $01e91
          7826 => x"81", -- $01e92
          7827 => x"80", -- $01e93
          7828 => x"7f", -- $01e94
          7829 => x"7e", -- $01e95
          7830 => x"7e", -- $01e96
          7831 => x"7d", -- $01e97
          7832 => x"7d", -- $01e98
          7833 => x"7e", -- $01e99
          7834 => x"7e", -- $01e9a
          7835 => x"7e", -- $01e9b
          7836 => x"7e", -- $01e9c
          7837 => x"7e", -- $01e9d
          7838 => x"7d", -- $01e9e
          7839 => x"7d", -- $01e9f
          7840 => x"7e", -- $01ea0
          7841 => x"7d", -- $01ea1
          7842 => x"7d", -- $01ea2
          7843 => x"7e", -- $01ea3
          7844 => x"7e", -- $01ea4
          7845 => x"7e", -- $01ea5
          7846 => x"7d", -- $01ea6
          7847 => x"7d", -- $01ea7
          7848 => x"7d", -- $01ea8
          7849 => x"7d", -- $01ea9
          7850 => x"7d", -- $01eaa
          7851 => x"7c", -- $01eab
          7852 => x"7c", -- $01eac
          7853 => x"7c", -- $01ead
          7854 => x"7c", -- $01eae
          7855 => x"7c", -- $01eaf
          7856 => x"7c", -- $01eb0
          7857 => x"7c", -- $01eb1
          7858 => x"7d", -- $01eb2
          7859 => x"7e", -- $01eb3
          7860 => x"7f", -- $01eb4
          7861 => x"80", -- $01eb5
          7862 => x"80", -- $01eb6
          7863 => x"81", -- $01eb7
          7864 => x"82", -- $01eb8
          7865 => x"82", -- $01eb9
          7866 => x"83", -- $01eba
          7867 => x"84", -- $01ebb
          7868 => x"84", -- $01ebc
          7869 => x"85", -- $01ebd
          7870 => x"86", -- $01ebe
          7871 => x"86", -- $01ebf
          7872 => x"87", -- $01ec0
          7873 => x"86", -- $01ec1
          7874 => x"85", -- $01ec2
          7875 => x"85", -- $01ec3
          7876 => x"84", -- $01ec4
          7877 => x"83", -- $01ec5
          7878 => x"82", -- $01ec6
          7879 => x"81", -- $01ec7
          7880 => x"82", -- $01ec8
          7881 => x"82", -- $01ec9
          7882 => x"83", -- $01eca
          7883 => x"83", -- $01ecb
          7884 => x"84", -- $01ecc
          7885 => x"85", -- $01ecd
          7886 => x"84", -- $01ece
          7887 => x"83", -- $01ecf
          7888 => x"81", -- $01ed0
          7889 => x"7f", -- $01ed1
          7890 => x"7d", -- $01ed2
          7891 => x"7b", -- $01ed3
          7892 => x"7b", -- $01ed4
          7893 => x"7b", -- $01ed5
          7894 => x"7d", -- $01ed6
          7895 => x"7e", -- $01ed7
          7896 => x"7f", -- $01ed8
          7897 => x"80", -- $01ed9
          7898 => x"7f", -- $01eda
          7899 => x"7d", -- $01edb
          7900 => x"7a", -- $01edc
          7901 => x"78", -- $01edd
          7902 => x"78", -- $01ede
          7903 => x"78", -- $01edf
          7904 => x"79", -- $01ee0
          7905 => x"7c", -- $01ee1
          7906 => x"7e", -- $01ee2
          7907 => x"80", -- $01ee3
          7908 => x"82", -- $01ee4
          7909 => x"82", -- $01ee5
          7910 => x"82", -- $01ee6
          7911 => x"81", -- $01ee7
          7912 => x"80", -- $01ee8
          7913 => x"80", -- $01ee9
          7914 => x"7f", -- $01eea
          7915 => x"7f", -- $01eeb
          7916 => x"7e", -- $01eec
          7917 => x"7e", -- $01eed
          7918 => x"7e", -- $01eee
          7919 => x"7d", -- $01eef
          7920 => x"7c", -- $01ef0
          7921 => x"7c", -- $01ef1
          7922 => x"7b", -- $01ef2
          7923 => x"7b", -- $01ef3
          7924 => x"7c", -- $01ef4
          7925 => x"7d", -- $01ef5
          7926 => x"7d", -- $01ef6
          7927 => x"7e", -- $01ef7
          7928 => x"7e", -- $01ef8
          7929 => x"7f", -- $01ef9
          7930 => x"80", -- $01efa
          7931 => x"80", -- $01efb
          7932 => x"80", -- $01efc
          7933 => x"80", -- $01efd
          7934 => x"80", -- $01efe
          7935 => x"80", -- $01eff
          7936 => x"80", -- $01f00
          7937 => x"80", -- $01f01
          7938 => x"80", -- $01f02
          7939 => x"81", -- $01f03
          7940 => x"82", -- $01f04
          7941 => x"83", -- $01f05
          7942 => x"84", -- $01f06
          7943 => x"84", -- $01f07
          7944 => x"85", -- $01f08
          7945 => x"85", -- $01f09
          7946 => x"86", -- $01f0a
          7947 => x"86", -- $01f0b
          7948 => x"87", -- $01f0c
          7949 => x"87", -- $01f0d
          7950 => x"86", -- $01f0e
          7951 => x"86", -- $01f0f
          7952 => x"85", -- $01f10
          7953 => x"85", -- $01f11
          7954 => x"84", -- $01f12
          7955 => x"84", -- $01f13
          7956 => x"84", -- $01f14
          7957 => x"83", -- $01f15
          7958 => x"82", -- $01f16
          7959 => x"80", -- $01f17
          7960 => x"7e", -- $01f18
          7961 => x"7c", -- $01f19
          7962 => x"7c", -- $01f1a
          7963 => x"7d", -- $01f1b
          7964 => x"7d", -- $01f1c
          7965 => x"7f", -- $01f1d
          7966 => x"7f", -- $01f1e
          7967 => x"7f", -- $01f1f
          7968 => x"7d", -- $01f20
          7969 => x"7a", -- $01f21
          7970 => x"77", -- $01f22
          7971 => x"75", -- $01f23
          7972 => x"74", -- $01f24
          7973 => x"75", -- $01f25
          7974 => x"77", -- $01f26
          7975 => x"79", -- $01f27
          7976 => x"7c", -- $01f28
          7977 => x"7e", -- $01f29
          7978 => x"7f", -- $01f2a
          7979 => x"7f", -- $01f2b
          7980 => x"7e", -- $01f2c
          7981 => x"7d", -- $01f2d
          7982 => x"7c", -- $01f2e
          7983 => x"7b", -- $01f2f
          7984 => x"7b", -- $01f30
          7985 => x"7b", -- $01f31
          7986 => x"7b", -- $01f32
          7987 => x"7c", -- $01f33
          7988 => x"7c", -- $01f34
          7989 => x"7c", -- $01f35
          7990 => x"7d", -- $01f36
          7991 => x"7e", -- $01f37
          7992 => x"7f", -- $01f38
          7993 => x"80", -- $01f39
          7994 => x"80", -- $01f3a
          7995 => x"81", -- $01f3b
          7996 => x"82", -- $01f3c
          7997 => x"82", -- $01f3d
          7998 => x"81", -- $01f3e
          7999 => x"81", -- $01f3f
          8000 => x"81", -- $01f40
          8001 => x"81", -- $01f41
          8002 => x"81", -- $01f42
          8003 => x"80", -- $01f43
          8004 => x"80", -- $01f44
          8005 => x"80", -- $01f45
          8006 => x"7f", -- $01f46
          8007 => x"7e", -- $01f47
          8008 => x"7e", -- $01f48
          8009 => x"7e", -- $01f49
          8010 => x"7f", -- $01f4a
          8011 => x"80", -- $01f4b
          8012 => x"80", -- $01f4c
          8013 => x"81", -- $01f4d
          8014 => x"83", -- $01f4e
          8015 => x"83", -- $01f4f
          8016 => x"84", -- $01f50
          8017 => x"85", -- $01f51
          8018 => x"85", -- $01f52
          8019 => x"85", -- $01f53
          8020 => x"86", -- $01f54
          8021 => x"86", -- $01f55
          8022 => x"86", -- $01f56
          8023 => x"84", -- $01f57
          8024 => x"84", -- $01f58
          8025 => x"81", -- $01f59
          8026 => x"80", -- $01f5a
          8027 => x"80", -- $01f5b
          8028 => x"80", -- $01f5c
          8029 => x"82", -- $01f5d
          8030 => x"82", -- $01f5e
          8031 => x"83", -- $01f5f
          8032 => x"82", -- $01f60
          8033 => x"80", -- $01f61
          8034 => x"7d", -- $01f62
          8035 => x"78", -- $01f63
          8036 => x"75", -- $01f64
          8037 => x"72", -- $01f65
          8038 => x"72", -- $01f66
          8039 => x"74", -- $01f67
          8040 => x"76", -- $01f68
          8041 => x"78", -- $01f69
          8042 => x"7a", -- $01f6a
          8043 => x"7c", -- $01f6b
          8044 => x"7c", -- $01f6c
          8045 => x"7c", -- $01f6d
          8046 => x"7c", -- $01f6e
          8047 => x"7b", -- $01f6f
          8048 => x"7b", -- $01f70
          8049 => x"7a", -- $01f71
          8050 => x"79", -- $01f72
          8051 => x"78", -- $01f73
          8052 => x"78", -- $01f74
          8053 => x"79", -- $01f75
          8054 => x"79", -- $01f76
          8055 => x"7a", -- $01f77
          8056 => x"7b", -- $01f78
          8057 => x"7c", -- $01f79
          8058 => x"7e", -- $01f7a
          8059 => x"7e", -- $01f7b
          8060 => x"7e", -- $01f7c
          8061 => x"7f", -- $01f7d
          8062 => x"80", -- $01f7e
          8063 => x"81", -- $01f7f
          8064 => x"83", -- $01f80
          8065 => x"84", -- $01f81
          8066 => x"86", -- $01f82
          8067 => x"86", -- $01f83
          8068 => x"85", -- $01f84
          8069 => x"84", -- $01f85
          8070 => x"83", -- $01f86
          8071 => x"81", -- $01f87
          8072 => x"80", -- $01f88
          8073 => x"80", -- $01f89
          8074 => x"80", -- $01f8a
          8075 => x"80", -- $01f8b
          8076 => x"7f", -- $01f8c
          8077 => x"80", -- $01f8d
          8078 => x"80", -- $01f8e
          8079 => x"80", -- $01f8f
          8080 => x"81", -- $01f90
          8081 => x"82", -- $01f91
          8082 => x"82", -- $01f92
          8083 => x"82", -- $01f93
          8084 => x"82", -- $01f94
          8085 => x"82", -- $01f95
          8086 => x"81", -- $01f96
          8087 => x"80", -- $01f97
          8088 => x"80", -- $01f98
          8089 => x"7f", -- $01f99
          8090 => x"7f", -- $01f9a
          8091 => x"80", -- $01f9b
          8092 => x"80", -- $01f9c
          8093 => x"81", -- $01f9d
          8094 => x"83", -- $01f9e
          8095 => x"83", -- $01f9f
          8096 => x"84", -- $01fa0
          8097 => x"82", -- $01fa1
          8098 => x"80", -- $01fa2
          8099 => x"7e", -- $01fa3
          8100 => x"7b", -- $01fa4
          8101 => x"7a", -- $01fa5
          8102 => x"78", -- $01fa6
          8103 => x"77", -- $01fa7
          8104 => x"78", -- $01fa8
          8105 => x"79", -- $01fa9
          8106 => x"7a", -- $01faa
          8107 => x"7c", -- $01fab
          8108 => x"7d", -- $01fac
          8109 => x"7e", -- $01fad
          8110 => x"7e", -- $01fae
          8111 => x"7f", -- $01faf
          8112 => x"7e", -- $01fb0
          8113 => x"7c", -- $01fb1
          8114 => x"7b", -- $01fb2
          8115 => x"79", -- $01fb3
          8116 => x"78", -- $01fb4
          8117 => x"79", -- $01fb5
          8118 => x"7a", -- $01fb6
          8119 => x"7b", -- $01fb7
          8120 => x"7d", -- $01fb8
          8121 => x"7e", -- $01fb9
          8122 => x"7e", -- $01fba
          8123 => x"7e", -- $01fbb
          8124 => x"7d", -- $01fbc
          8125 => x"7d", -- $01fbd
          8126 => x"7d", -- $01fbe
          8127 => x"7e", -- $01fbf
          8128 => x"80", -- $01fc0
          8129 => x"82", -- $01fc1
          8130 => x"84", -- $01fc2
          8131 => x"85", -- $01fc3
          8132 => x"85", -- $01fc4
          8133 => x"86", -- $01fc5
          8134 => x"85", -- $01fc6
          8135 => x"84", -- $01fc7
          8136 => x"84", -- $01fc8
          8137 => x"82", -- $01fc9
          8138 => x"82", -- $01fca
          8139 => x"81", -- $01fcb
          8140 => x"81", -- $01fcc
          8141 => x"82", -- $01fcd
          8142 => x"83", -- $01fce
          8143 => x"86", -- $01fcf
          8144 => x"87", -- $01fd0
          8145 => x"88", -- $01fd1
          8146 => x"87", -- $01fd2
          8147 => x"86", -- $01fd3
          8148 => x"86", -- $01fd4
          8149 => x"85", -- $01fd5
          8150 => x"86", -- $01fd6
          8151 => x"84", -- $01fd7
          8152 => x"84", -- $01fd8
          8153 => x"82", -- $01fd9
          8154 => x"80", -- $01fda
          8155 => x"80", -- $01fdb
          8156 => x"80", -- $01fdc
          8157 => x"82", -- $01fdd
          8158 => x"83", -- $01fde
          8159 => x"85", -- $01fdf
          8160 => x"84", -- $01fe0
          8161 => x"82", -- $01fe1
          8162 => x"7e", -- $01fe2
          8163 => x"79", -- $01fe3
          8164 => x"75", -- $01fe4
          8165 => x"72", -- $01fe5
          8166 => x"72", -- $01fe6
          8167 => x"73", -- $01fe7
          8168 => x"76", -- $01fe8
          8169 => x"79", -- $01fe9
          8170 => x"7b", -- $01fea
          8171 => x"7e", -- $01feb
          8172 => x"7f", -- $01fec
          8173 => x"7f", -- $01fed
          8174 => x"7f", -- $01fee
          8175 => x"7d", -- $01fef
          8176 => x"7c", -- $01ff0
          8177 => x"7b", -- $01ff1
          8178 => x"7a", -- $01ff2
          8179 => x"7a", -- $01ff3
          8180 => x"7b", -- $01ff4
          8181 => x"7e", -- $01ff5
          8182 => x"80", -- $01ff6
          8183 => x"81", -- $01ff7
          8184 => x"81", -- $01ff8
          8185 => x"81", -- $01ff9
          8186 => x"80", -- $01ffa
          8187 => x"7f", -- $01ffb
          8188 => x"7f", -- $01ffc
          8189 => x"7f", -- $01ffd
          8190 => x"80", -- $01ffe
          8191 => x"81", -- $01fff
          8192 => x"83", -- $02000
          8193 => x"83", -- $02001
          8194 => x"83", -- $02002
          8195 => x"84", -- $02003
          8196 => x"83", -- $02004
          8197 => x"84", -- $02005
          8198 => x"82", -- $02006
          8199 => x"82", -- $02007
          8200 => x"82", -- $02008
          8201 => x"81", -- $02009
          8202 => x"83", -- $0200a
          8203 => x"83", -- $0200b
          8204 => x"84", -- $0200c
          8205 => x"84", -- $0200d
          8206 => x"85", -- $0200e
          8207 => x"85", -- $0200f
          8208 => x"85", -- $02010
          8209 => x"86", -- $02011
          8210 => x"86", -- $02012
          8211 => x"86", -- $02013
          8212 => x"86", -- $02014
          8213 => x"83", -- $02015
          8214 => x"83", -- $02016
          8215 => x"81", -- $02017
          8216 => x"82", -- $02018
          8217 => x"84", -- $02019
          8218 => x"86", -- $0201a
          8219 => x"88", -- $0201b
          8220 => x"87", -- $0201c
          8221 => x"84", -- $0201d
          8222 => x"80", -- $0201e
          8223 => x"7b", -- $0201f
          8224 => x"77", -- $02020
          8225 => x"74", -- $02021
          8226 => x"75", -- $02022
          8227 => x"76", -- $02023
          8228 => x"78", -- $02024
          8229 => x"7a", -- $02025
          8230 => x"7c", -- $02026
          8231 => x"7d", -- $02027
          8232 => x"7e", -- $02028
          8233 => x"7e", -- $02029
          8234 => x"7d", -- $0202a
          8235 => x"7c", -- $0202b
          8236 => x"7a", -- $0202c
          8237 => x"79", -- $0202d
          8238 => x"78", -- $0202e
          8239 => x"79", -- $0202f
          8240 => x"7a", -- $02030
          8241 => x"7c", -- $02031
          8242 => x"7e", -- $02032
          8243 => x"80", -- $02033
          8244 => x"80", -- $02034
          8245 => x"7f", -- $02035
          8246 => x"7f", -- $02036
          8247 => x"7e", -- $02037
          8248 => x"7f", -- $02038
          8249 => x"80", -- $02039
          8250 => x"81", -- $0203a
          8251 => x"82", -- $0203b
          8252 => x"83", -- $0203c
          8253 => x"84", -- $0203d
          8254 => x"84", -- $0203e
          8255 => x"83", -- $0203f
          8256 => x"83", -- $02040
          8257 => x"83", -- $02041
          8258 => x"83", -- $02042
          8259 => x"84", -- $02043
          8260 => x"84", -- $02044
          8261 => x"85", -- $02045
          8262 => x"85", -- $02046
          8263 => x"85", -- $02047
          8264 => x"85", -- $02048
          8265 => x"84", -- $02049
          8266 => x"85", -- $0204a
          8267 => x"86", -- $0204b
          8268 => x"86", -- $0204c
          8269 => x"87", -- $0204d
          8270 => x"85", -- $0204e
          8271 => x"85", -- $0204f
          8272 => x"82", -- $02050
          8273 => x"80", -- $02051
          8274 => x"81", -- $02052
          8275 => x"81", -- $02053
          8276 => x"84", -- $02054
          8277 => x"87", -- $02055
          8278 => x"89", -- $02056
          8279 => x"88", -- $02057
          8280 => x"84", -- $02058
          8281 => x"80", -- $02059
          8282 => x"7b", -- $0205a
          8283 => x"77", -- $0205b
          8284 => x"75", -- $0205c
          8285 => x"74", -- $0205d
          8286 => x"76", -- $0205e
          8287 => x"78", -- $0205f
          8288 => x"7b", -- $02060
          8289 => x"7d", -- $02061
          8290 => x"7f", -- $02062
          8291 => x"80", -- $02063
          8292 => x"7f", -- $02064
          8293 => x"7f", -- $02065
          8294 => x"7c", -- $02066
          8295 => x"7b", -- $02067
          8296 => x"7a", -- $02068
          8297 => x"7a", -- $02069
          8298 => x"7c", -- $0206a
          8299 => x"7e", -- $0206b
          8300 => x"80", -- $0206c
          8301 => x"80", -- $0206d
          8302 => x"81", -- $0206e
          8303 => x"81", -- $0206f
          8304 => x"80", -- $02070
          8305 => x"80", -- $02071
          8306 => x"7f", -- $02072
          8307 => x"7f", -- $02073
          8308 => x"80", -- $02074
          8309 => x"80", -- $02075
          8310 => x"81", -- $02076
          8311 => x"82", -- $02077
          8312 => x"83", -- $02078
          8313 => x"84", -- $02079
          8314 => x"85", -- $0207a
          8315 => x"84", -- $0207b
          8316 => x"83", -- $0207c
          8317 => x"83", -- $0207d
          8318 => x"82", -- $0207e
          8319 => x"82", -- $0207f
          8320 => x"82", -- $02080
          8321 => x"82", -- $02081
          8322 => x"81", -- $02082
          8323 => x"82", -- $02083
          8324 => x"82", -- $02084
          8325 => x"84", -- $02085
          8326 => x"87", -- $02086
          8327 => x"87", -- $02087
          8328 => x"85", -- $02088
          8329 => x"83", -- $02089
          8330 => x"81", -- $0208a
          8331 => x"81", -- $0208b
          8332 => x"83", -- $0208c
          8333 => x"87", -- $0208d
          8334 => x"8b", -- $0208e
          8335 => x"8d", -- $0208f
          8336 => x"8d", -- $02090
          8337 => x"89", -- $02091
          8338 => x"84", -- $02092
          8339 => x"7f", -- $02093
          8340 => x"7b", -- $02094
          8341 => x"79", -- $02095
          8342 => x"7a", -- $02096
          8343 => x"7c", -- $02097
          8344 => x"7d", -- $02098
          8345 => x"7e", -- $02099
          8346 => x"7e", -- $0209a
          8347 => x"7e", -- $0209b
          8348 => x"7e", -- $0209c
          8349 => x"7d", -- $0209d
          8350 => x"7c", -- $0209e
          8351 => x"7b", -- $0209f
          8352 => x"7b", -- $020a0
          8353 => x"7b", -- $020a1
          8354 => x"7c", -- $020a2
          8355 => x"7d", -- $020a3
          8356 => x"7f", -- $020a4
          8357 => x"81", -- $020a5
          8358 => x"82", -- $020a6
          8359 => x"82", -- $020a7
          8360 => x"81", -- $020a8
          8361 => x"80", -- $020a9
          8362 => x"80", -- $020aa
          8363 => x"80", -- $020ab
          8364 => x"81", -- $020ac
          8365 => x"82", -- $020ad
          8366 => x"82", -- $020ae
          8367 => x"82", -- $020af
          8368 => x"83", -- $020b0
          8369 => x"83", -- $020b1
          8370 => x"82", -- $020b2
          8371 => x"82", -- $020b3
          8372 => x"82", -- $020b4
          8373 => x"82", -- $020b5
          8374 => x"82", -- $020b6
          8375 => x"82", -- $020b7
          8376 => x"83", -- $020b8
          8377 => x"83", -- $020b9
          8378 => x"85", -- $020ba
          8379 => x"86", -- $020bb
          8380 => x"88", -- $020bc
          8381 => x"85", -- $020bd
          8382 => x"81", -- $020be
          8383 => x"80", -- $020bf
          8384 => x"7e", -- $020c0
          8385 => x"80", -- $020c1
          8386 => x"83", -- $020c2
          8387 => x"86", -- $020c3
          8388 => x"8a", -- $020c4
          8389 => x"8a", -- $020c5
          8390 => x"88", -- $020c6
          8391 => x"83", -- $020c7
          8392 => x"7f", -- $020c8
          8393 => x"7c", -- $020c9
          8394 => x"7a", -- $020ca
          8395 => x"7b", -- $020cb
          8396 => x"7d", -- $020cc
          8397 => x"7f", -- $020cd
          8398 => x"80", -- $020ce
          8399 => x"80", -- $020cf
          8400 => x"80", -- $020d0
          8401 => x"81", -- $020d1
          8402 => x"80", -- $020d2
          8403 => x"80", -- $020d3
          8404 => x"80", -- $020d4
          8405 => x"7f", -- $020d5
          8406 => x"7e", -- $020d6
          8407 => x"7e", -- $020d7
          8408 => x"7f", -- $020d8
          8409 => x"80", -- $020d9
          8410 => x"82", -- $020da
          8411 => x"83", -- $020db
          8412 => x"84", -- $020dc
          8413 => x"84", -- $020dd
          8414 => x"82", -- $020de
          8415 => x"81", -- $020df
          8416 => x"80", -- $020e0
          8417 => x"80", -- $020e1
          8418 => x"80", -- $020e2
          8419 => x"80", -- $020e3
          8420 => x"80", -- $020e4
          8421 => x"80", -- $020e5
          8422 => x"80", -- $020e6
          8423 => x"80", -- $020e7
          8424 => x"80", -- $020e8
          8425 => x"7f", -- $020e9
          8426 => x"7e", -- $020ea
          8427 => x"7e", -- $020eb
          8428 => x"7e", -- $020ec
          8429 => x"7f", -- $020ed
          8430 => x"7f", -- $020ee
          8431 => x"80", -- $020ef
          8432 => x"81", -- $020f0
          8433 => x"84", -- $020f1
          8434 => x"84", -- $020f2
          8435 => x"7f", -- $020f3
          8436 => x"7e", -- $020f4
          8437 => x"7d", -- $020f5
          8438 => x"7c", -- $020f6
          8439 => x"80", -- $020f7
          8440 => x"83", -- $020f8
          8441 => x"88", -- $020f9
          8442 => x"89", -- $020fa
          8443 => x"86", -- $020fb
          8444 => x"85", -- $020fc
          8445 => x"80", -- $020fd
          8446 => x"7b", -- $020fe
          8447 => x"7a", -- $020ff
          8448 => x"7b", -- $02100
          8449 => x"7c", -- $02101
          8450 => x"80", -- $02102
          8451 => x"81", -- $02103
          8452 => x"82", -- $02104
          8453 => x"81", -- $02105
          8454 => x"82", -- $02106
          8455 => x"83", -- $02107
          8456 => x"81", -- $02108
          8457 => x"81", -- $02109
          8458 => x"81", -- $0210a
          8459 => x"80", -- $0210b
          8460 => x"80", -- $0210c
          8461 => x"80", -- $0210d
          8462 => x"82", -- $0210e
          8463 => x"83", -- $0210f
          8464 => x"84", -- $02110
          8465 => x"86", -- $02111
          8466 => x"86", -- $02112
          8467 => x"84", -- $02113
          8468 => x"83", -- $02114
          8469 => x"82", -- $02115
          8470 => x"81", -- $02116
          8471 => x"81", -- $02117
          8472 => x"82", -- $02118
          8473 => x"82", -- $02119
          8474 => x"83", -- $0211a
          8475 => x"82", -- $0211b
          8476 => x"81", -- $0211c
          8477 => x"81", -- $0211d
          8478 => x"80", -- $0211e
          8479 => x"7f", -- $0211f
          8480 => x"7f", -- $02120
          8481 => x"7f", -- $02121
          8482 => x"80", -- $02122
          8483 => x"7f", -- $02123
          8484 => x"80", -- $02124
          8485 => x"81", -- $02125
          8486 => x"80", -- $02126
          8487 => x"7e", -- $02127
          8488 => x"7d", -- $02128
          8489 => x"7d", -- $02129
          8490 => x"7d", -- $0212a
          8491 => x"7f", -- $0212b
          8492 => x"80", -- $0212c
          8493 => x"83", -- $0212d
          8494 => x"84", -- $0212e
          8495 => x"82", -- $0212f
          8496 => x"80", -- $02130
          8497 => x"7e", -- $02131
          8498 => x"7b", -- $02132
          8499 => x"79", -- $02133
          8500 => x"7a", -- $02134
          8501 => x"7c", -- $02135
          8502 => x"7f", -- $02136
          8503 => x"80", -- $02137
          8504 => x"81", -- $02138
          8505 => x"82", -- $02139
          8506 => x"81", -- $0213a
          8507 => x"81", -- $0213b
          8508 => x"80", -- $0213c
          8509 => x"80", -- $0213d
          8510 => x"80", -- $0213e
          8511 => x"80", -- $0213f
          8512 => x"81", -- $02140
          8513 => x"82", -- $02141
          8514 => x"83", -- $02142
          8515 => x"84", -- $02143
          8516 => x"84", -- $02144
          8517 => x"85", -- $02145
          8518 => x"86", -- $02146
          8519 => x"85", -- $02147
          8520 => x"84", -- $02148
          8521 => x"84", -- $02149
          8522 => x"84", -- $0214a
          8523 => x"84", -- $0214b
          8524 => x"84", -- $0214c
          8525 => x"84", -- $0214d
          8526 => x"85", -- $0214e
          8527 => x"85", -- $0214f
          8528 => x"85", -- $02150
          8529 => x"84", -- $02151
          8530 => x"83", -- $02152
          8531 => x"82", -- $02153
          8532 => x"81", -- $02154
          8533 => x"80", -- $02155
          8534 => x"80", -- $02156
          8535 => x"7f", -- $02157
          8536 => x"7f", -- $02158
          8537 => x"7f", -- $02159
          8538 => x"7e", -- $0215a
          8539 => x"7e", -- $0215b
          8540 => x"7e", -- $0215c
          8541 => x"7e", -- $0215d
          8542 => x"7e", -- $0215e
          8543 => x"7d", -- $0215f
          8544 => x"7d", -- $02160
          8545 => x"7d", -- $02161
          8546 => x"7c", -- $02162
          8547 => x"7b", -- $02163
          8548 => x"7a", -- $02164
          8549 => x"79", -- $02165
          8550 => x"79", -- $02166
          8551 => x"79", -- $02167
          8552 => x"7a", -- $02168
          8553 => x"7a", -- $02169
          8554 => x"7c", -- $0216a
          8555 => x"7c", -- $0216b
          8556 => x"7d", -- $0216c
          8557 => x"7e", -- $0216d
          8558 => x"7e", -- $0216e
          8559 => x"7f", -- $0216f
          8560 => x"80", -- $02170
          8561 => x"80", -- $02171
          8562 => x"81", -- $02172
          8563 => x"82", -- $02173
          8564 => x"83", -- $02174
          8565 => x"85", -- $02175
          8566 => x"87", -- $02176
          8567 => x"8a", -- $02177
          8568 => x"8c", -- $02178
          8569 => x"8e", -- $02179
          8570 => x"8f", -- $0217a
          8571 => x"8e", -- $0217b
          8572 => x"8c", -- $0217c
          8573 => x"89", -- $0217d
          8574 => x"87", -- $0217e
          8575 => x"86", -- $0217f
          8576 => x"87", -- $02180
          8577 => x"88", -- $02181
          8578 => x"89", -- $02182
          8579 => x"88", -- $02183
          8580 => x"86", -- $02184
          8581 => x"84", -- $02185
          8582 => x"80", -- $02186
          8583 => x"7c", -- $02187
          8584 => x"78", -- $02188
          8585 => x"76", -- $02189
          8586 => x"75", -- $0218a
          8587 => x"75", -- $0218b
          8588 => x"75", -- $0218c
          8589 => x"75", -- $0218d
          8590 => x"75", -- $0218e
          8591 => x"76", -- $0218f
          8592 => x"77", -- $02190
          8593 => x"78", -- $02191
          8594 => x"7a", -- $02192
          8595 => x"7c", -- $02193
          8596 => x"7e", -- $02194
          8597 => x"80", -- $02195
          8598 => x"80", -- $02196
          8599 => x"81", -- $02197
          8600 => x"81", -- $02198
          8601 => x"81", -- $02199
          8602 => x"81", -- $0219a
          8603 => x"81", -- $0219b
          8604 => x"80", -- $0219c
          8605 => x"80", -- $0219d
          8606 => x"7f", -- $0219e
          8607 => x"7e", -- $0219f
          8608 => x"7f", -- $021a0
          8609 => x"7f", -- $021a1
          8610 => x"7f", -- $021a2
          8611 => x"80", -- $021a3
          8612 => x"80", -- $021a4
          8613 => x"80", -- $021a5
          8614 => x"80", -- $021a6
          8615 => x"81", -- $021a7
          8616 => x"82", -- $021a8
          8617 => x"83", -- $021a9
          8618 => x"84", -- $021aa
          8619 => x"85", -- $021ab
          8620 => x"85", -- $021ac
          8621 => x"85", -- $021ad
          8622 => x"84", -- $021ae
          8623 => x"83", -- $021af
          8624 => x"82", -- $021b0
          8625 => x"81", -- $021b1
          8626 => x"80", -- $021b2
          8627 => x"80", -- $021b3
          8628 => x"81", -- $021b4
          8629 => x"81", -- $021b5
          8630 => x"82", -- $021b6
          8631 => x"82", -- $021b7
          8632 => x"82", -- $021b8
          8633 => x"81", -- $021b9
          8634 => x"81", -- $021ba
          8635 => x"80", -- $021bb
          8636 => x"80", -- $021bc
          8637 => x"80", -- $021bd
          8638 => x"80", -- $021be
          8639 => x"7f", -- $021bf
          8640 => x"7f", -- $021c0
          8641 => x"7e", -- $021c1
          8642 => x"7e", -- $021c2
          8643 => x"7d", -- $021c3
          8644 => x"7d", -- $021c4
          8645 => x"7c", -- $021c5
          8646 => x"7c", -- $021c6
          8647 => x"7c", -- $021c7
          8648 => x"7b", -- $021c8
          8649 => x"7b", -- $021c9
          8650 => x"7b", -- $021ca
          8651 => x"7c", -- $021cb
          8652 => x"7c", -- $021cc
          8653 => x"7d", -- $021cd
          8654 => x"7f", -- $021ce
          8655 => x"80", -- $021cf
          8656 => x"80", -- $021d0
          8657 => x"81", -- $021d1
          8658 => x"82", -- $021d2
          8659 => x"83", -- $021d3
          8660 => x"84", -- $021d4
          8661 => x"86", -- $021d5
          8662 => x"88", -- $021d6
          8663 => x"89", -- $021d7
          8664 => x"89", -- $021d8
          8665 => x"86", -- $021d9
          8666 => x"84", -- $021da
          8667 => x"82", -- $021db
          8668 => x"80", -- $021dc
          8669 => x"80", -- $021dd
          8670 => x"81", -- $021de
          8671 => x"83", -- $021df
          8672 => x"84", -- $021e0
          8673 => x"83", -- $021e1
          8674 => x"82", -- $021e2
          8675 => x"80", -- $021e3
          8676 => x"7c", -- $021e4
          8677 => x"79", -- $021e5
          8678 => x"77", -- $021e6
          8679 => x"77", -- $021e7
          8680 => x"78", -- $021e8
          8681 => x"78", -- $021e9
          8682 => x"79", -- $021ea
          8683 => x"7a", -- $021eb
          8684 => x"7a", -- $021ec
          8685 => x"7a", -- $021ed
          8686 => x"7b", -- $021ee
          8687 => x"7d", -- $021ef
          8688 => x"7e", -- $021f0
          8689 => x"7f", -- $021f1
          8690 => x"80", -- $021f2
          8691 => x"81", -- $021f3
          8692 => x"82", -- $021f4
          8693 => x"82", -- $021f5
          8694 => x"82", -- $021f6
          8695 => x"82", -- $021f7
          8696 => x"82", -- $021f8
          8697 => x"81", -- $021f9
          8698 => x"80", -- $021fa
          8699 => x"80", -- $021fb
          8700 => x"80", -- $021fc
          8701 => x"7f", -- $021fd
          8702 => x"7f", -- $021fe
          8703 => x"7f", -- $021ff
          8704 => x"80", -- $02200
          8705 => x"80", -- $02201
          8706 => x"80", -- $02202
          8707 => x"80", -- $02203
          8708 => x"81", -- $02204
          8709 => x"81", -- $02205
          8710 => x"81", -- $02206
          8711 => x"81", -- $02207
          8712 => x"81", -- $02208
          8713 => x"80", -- $02209
          8714 => x"80", -- $0220a
          8715 => x"7f", -- $0220b
          8716 => x"7e", -- $0220c
          8717 => x"7e", -- $0220d
          8718 => x"7e", -- $0220e
          8719 => x"7f", -- $0220f
          8720 => x"80", -- $02210
          8721 => x"80", -- $02211
          8722 => x"80", -- $02212
          8723 => x"80", -- $02213
          8724 => x"80", -- $02214
          8725 => x"80", -- $02215
          8726 => x"80", -- $02216
          8727 => x"80", -- $02217
          8728 => x"80", -- $02218
          8729 => x"80", -- $02219
          8730 => x"80", -- $0221a
          8731 => x"7f", -- $0221b
          8732 => x"7e", -- $0221c
          8733 => x"7c", -- $0221d
          8734 => x"7b", -- $0221e
          8735 => x"7b", -- $0221f
          8736 => x"7a", -- $02220
          8737 => x"79", -- $02221
          8738 => x"78", -- $02222
          8739 => x"77", -- $02223
          8740 => x"76", -- $02224
          8741 => x"75", -- $02225
          8742 => x"75", -- $02226
          8743 => x"76", -- $02227
          8744 => x"78", -- $02228
          8745 => x"7a", -- $02229
          8746 => x"7d", -- $0222a
          8747 => x"7e", -- $0222b
          8748 => x"80", -- $0222c
          8749 => x"82", -- $0222d
          8750 => x"85", -- $0222e
          8751 => x"87", -- $0222f
          8752 => x"88", -- $02230
          8753 => x"8b", -- $02231
          8754 => x"8d", -- $02232
          8755 => x"8d", -- $02233
          8756 => x"8b", -- $02234
          8757 => x"89", -- $02235
          8758 => x"87", -- $02236
          8759 => x"83", -- $02237
          8760 => x"82", -- $02238
          8761 => x"83", -- $02239
          8762 => x"83", -- $0223a
          8763 => x"84", -- $0223b
          8764 => x"84", -- $0223c
          8765 => x"82", -- $0223d
          8766 => x"80", -- $0223e
          8767 => x"7b", -- $0223f
          8768 => x"77", -- $02240
          8769 => x"75", -- $02241
          8770 => x"73", -- $02242
          8771 => x"74", -- $02243
          8772 => x"77", -- $02244
          8773 => x"79", -- $02245
          8774 => x"7a", -- $02246
          8775 => x"7b", -- $02247
          8776 => x"7c", -- $02248
          8777 => x"7d", -- $02249
          8778 => x"7e", -- $0224a
          8779 => x"7f", -- $0224b
          8780 => x"80", -- $0224c
          8781 => x"80", -- $0224d
          8782 => x"81", -- $0224e
          8783 => x"81", -- $0224f
          8784 => x"81", -- $02250
          8785 => x"80", -- $02251
          8786 => x"80", -- $02252
          8787 => x"7f", -- $02253
          8788 => x"7f", -- $02254
          8789 => x"7e", -- $02255
          8790 => x"7d", -- $02256
          8791 => x"7d", -- $02257
          8792 => x"7c", -- $02258
          8793 => x"7b", -- $02259
          8794 => x"7c", -- $0225a
          8795 => x"7d", -- $0225b
          8796 => x"7e", -- $0225c
          8797 => x"80", -- $0225d
          8798 => x"80", -- $0225e
          8799 => x"80", -- $0225f
          8800 => x"81", -- $02260
          8801 => x"82", -- $02261
          8802 => x"84", -- $02262
          8803 => x"84", -- $02263
          8804 => x"84", -- $02264
          8805 => x"85", -- $02265
          8806 => x"83", -- $02266
          8807 => x"81", -- $02267
          8808 => x"81", -- $02268
          8809 => x"81", -- $02269
          8810 => x"81", -- $0226a
          8811 => x"81", -- $0226b
          8812 => x"84", -- $0226c
          8813 => x"84", -- $0226d
          8814 => x"84", -- $0226e
          8815 => x"83", -- $0226f
          8816 => x"83", -- $02270
          8817 => x"81", -- $02271
          8818 => x"80", -- $02272
          8819 => x"80", -- $02273
          8820 => x"80", -- $02274
          8821 => x"80", -- $02275
          8822 => x"80", -- $02276
          8823 => x"80", -- $02277
          8824 => x"80", -- $02278
          8825 => x"7e", -- $02279
          8826 => x"7d", -- $0227a
          8827 => x"7c", -- $0227b
          8828 => x"7b", -- $0227c
          8829 => x"7b", -- $0227d
          8830 => x"7b", -- $0227e
          8831 => x"7a", -- $0227f
          8832 => x"79", -- $02280
          8833 => x"79", -- $02281
          8834 => x"79", -- $02282
          8835 => x"7a", -- $02283
          8836 => x"7b", -- $02284
          8837 => x"7e", -- $02285
          8838 => x"7f", -- $02286
          8839 => x"80", -- $02287
          8840 => x"82", -- $02288
          8841 => x"83", -- $02289
          8842 => x"84", -- $0228a
          8843 => x"87", -- $0228b
          8844 => x"89", -- $0228c
          8845 => x"8c", -- $0228d
          8846 => x"8e", -- $0228e
          8847 => x"8f", -- $0228f
          8848 => x"8e", -- $02290
          8849 => x"86", -- $02291
          8850 => x"82", -- $02292
          8851 => x"7e", -- $02293
          8852 => x"7c", -- $02294
          8853 => x"7f", -- $02295
          8854 => x"82", -- $02296
          8855 => x"87", -- $02297
          8856 => x"88", -- $02298
          8857 => x"86", -- $02299
          8858 => x"81", -- $0229a
          8859 => x"7b", -- $0229b
          8860 => x"75", -- $0229c
          8861 => x"73", -- $0229d
          8862 => x"73", -- $0229e
          8863 => x"74", -- $0229f
          8864 => x"77", -- $022a0
          8865 => x"79", -- $022a1
          8866 => x"79", -- $022a2
          8867 => x"7a", -- $022a3
          8868 => x"7b", -- $022a4
          8869 => x"7d", -- $022a5
          8870 => x"80", -- $022a6
          8871 => x"82", -- $022a7
          8872 => x"84", -- $022a8
          8873 => x"81", -- $022a9
          8874 => x"80", -- $022aa
          8875 => x"7f", -- $022ab
          8876 => x"7e", -- $022ac
          8877 => x"7f", -- $022ad
          8878 => x"80", -- $022ae
          8879 => x"81", -- $022af
          8880 => x"81", -- $022b0
          8881 => x"80", -- $022b1
          8882 => x"7e", -- $022b2
          8883 => x"7d", -- $022b3
          8884 => x"7c", -- $022b4
          8885 => x"7d", -- $022b5
          8886 => x"7f", -- $022b6
          8887 => x"80", -- $022b7
          8888 => x"80", -- $022b8
          8889 => x"80", -- $022b9
          8890 => x"7f", -- $022ba
          8891 => x"7e", -- $022bb
          8892 => x"7f", -- $022bc
          8893 => x"80", -- $022bd
          8894 => x"82", -- $022be
          8895 => x"83", -- $022bf
          8896 => x"83", -- $022c0
          8897 => x"80", -- $022c1
          8898 => x"7e", -- $022c2
          8899 => x"7c", -- $022c3
          8900 => x"7c", -- $022c4
          8901 => x"7d", -- $022c5
          8902 => x"80", -- $022c6
          8903 => x"82", -- $022c7
          8904 => x"83", -- $022c8
          8905 => x"84", -- $022c9
          8906 => x"83", -- $022ca
          8907 => x"82", -- $022cb
          8908 => x"81", -- $022cc
          8909 => x"80", -- $022cd
          8910 => x"81", -- $022ce
          8911 => x"82", -- $022cf
          8912 => x"81", -- $022d0
          8913 => x"81", -- $022d1
          8914 => x"81", -- $022d2
          8915 => x"80", -- $022d3
          8916 => x"80", -- $022d4
          8917 => x"7e", -- $022d5
          8918 => x"7e", -- $022d6
          8919 => x"7d", -- $022d7
          8920 => x"7c", -- $022d8
          8921 => x"7b", -- $022d9
          8922 => x"7a", -- $022da
          8923 => x"79", -- $022db
          8924 => x"78", -- $022dc
          8925 => x"78", -- $022dd
          8926 => x"78", -- $022de
          8927 => x"77", -- $022df
          8928 => x"78", -- $022e0
          8929 => x"79", -- $022e1
          8930 => x"7a", -- $022e2
          8931 => x"7d", -- $022e3
          8932 => x"80", -- $022e4
          8933 => x"82", -- $022e5
          8934 => x"84", -- $022e6
          8935 => x"86", -- $022e7
          8936 => x"86", -- $022e8
          8937 => x"86", -- $022e9
          8938 => x"86", -- $022ea
          8939 => x"86", -- $022eb
          8940 => x"86", -- $022ec
          8941 => x"87", -- $022ed
          8942 => x"8a", -- $022ee
          8943 => x"8d", -- $022ef
          8944 => x"8e", -- $022f0
          8945 => x"8e", -- $022f1
          8946 => x"8a", -- $022f2
          8947 => x"7f", -- $022f3
          8948 => x"7a", -- $022f4
          8949 => x"77", -- $022f5
          8950 => x"76", -- $022f6
          8951 => x"7f", -- $022f7
          8952 => x"84", -- $022f8
          8953 => x"8a", -- $022f9
          8954 => x"8c", -- $022fa
          8955 => x"86", -- $022fb
          8956 => x"83", -- $022fc
          8957 => x"7e", -- $022fd
          8958 => x"7b", -- $022fe
          8959 => x"7c", -- $022ff
          8960 => x"7b", -- $02300
          8961 => x"7c", -- $02301
          8962 => x"79", -- $02302
          8963 => x"77", -- $02303
          8964 => x"77", -- $02304
          8965 => x"77", -- $02305
          8966 => x"7c", -- $02306
          8967 => x"82", -- $02307
          8968 => x"83", -- $02308
          8969 => x"85", -- $02309
          8970 => x"83", -- $0230a
          8971 => x"7f", -- $0230b
          8972 => x"7f", -- $0230c
          8973 => x"7e", -- $0230d
          8974 => x"7f", -- $0230e
          8975 => x"80", -- $0230f
          8976 => x"80", -- $02310
          8977 => x"7e", -- $02311
          8978 => x"7c", -- $02312
          8979 => x"7a", -- $02313
          8980 => x"7b", -- $02314
          8981 => x"7e", -- $02315
          8982 => x"80", -- $02316
          8983 => x"81", -- $02317
          8984 => x"81", -- $02318
          8985 => x"80", -- $02319
          8986 => x"7e", -- $0231a
          8987 => x"7e", -- $0231b
          8988 => x"80", -- $0231c
          8989 => x"81", -- $0231d
          8990 => x"84", -- $0231e
          8991 => x"86", -- $0231f
          8992 => x"86", -- $02320
          8993 => x"84", -- $02321
          8994 => x"84", -- $02322
          8995 => x"83", -- $02323
          8996 => x"83", -- $02324
          8997 => x"85", -- $02325
          8998 => x"85", -- $02326
          8999 => x"87", -- $02327
          9000 => x"87", -- $02328
          9001 => x"87", -- $02329
          9002 => x"8a", -- $0232a
          9003 => x"88", -- $0232b
          9004 => x"83", -- $0232c
          9005 => x"83", -- $0232d
          9006 => x"80", -- $0232e
          9007 => x"80", -- $0232f
          9008 => x"82", -- $02330
          9009 => x"84", -- $02331
          9010 => x"86", -- $02332
          9011 => x"85", -- $02333
          9012 => x"83", -- $02334
          9013 => x"80", -- $02335
          9014 => x"7e", -- $02336
          9015 => x"7d", -- $02337
          9016 => x"7a", -- $02338
          9017 => x"7a", -- $02339
          9018 => x"79", -- $0233a
          9019 => x"76", -- $0233b
          9020 => x"77", -- $0233c
          9021 => x"77", -- $0233d
          9022 => x"7b", -- $0233e
          9023 => x"7e", -- $0233f
          9024 => x"80", -- $02340
          9025 => x"80", -- $02341
          9026 => x"7d", -- $02342
          9027 => x"7b", -- $02343
          9028 => x"79", -- $02344
          9029 => x"7a", -- $02345
          9030 => x"7e", -- $02346
          9031 => x"80", -- $02347
          9032 => x"83", -- $02348
          9033 => x"83", -- $02349
          9034 => x"82", -- $0234a
          9035 => x"81", -- $0234b
          9036 => x"81", -- $0234c
          9037 => x"82", -- $0234d
          9038 => x"84", -- $0234e
          9039 => x"86", -- $0234f
          9040 => x"85", -- $02350
          9041 => x"83", -- $02351
          9042 => x"82", -- $02352
          9043 => x"82", -- $02353
          9044 => x"82", -- $02354
          9045 => x"83", -- $02355
          9046 => x"85", -- $02356
          9047 => x"84", -- $02357
          9048 => x"83", -- $02358
          9049 => x"82", -- $02359
          9050 => x"82", -- $0235a
          9051 => x"82", -- $0235b
          9052 => x"84", -- $0235c
          9053 => x"87", -- $0235d
          9054 => x"89", -- $0235e
          9055 => x"86", -- $0235f
          9056 => x"81", -- $02360
          9057 => x"80", -- $02361
          9058 => x"7c", -- $02362
          9059 => x"7f", -- $02363
          9060 => x"82", -- $02364
          9061 => x"86", -- $02365
          9062 => x"88", -- $02366
          9063 => x"85", -- $02367
          9064 => x"81", -- $02368
          9065 => x"7d", -- $02369
          9066 => x"7b", -- $0236a
          9067 => x"7b", -- $0236b
          9068 => x"7c", -- $0236c
          9069 => x"7d", -- $0236d
          9070 => x"7d", -- $0236e
          9071 => x"7b", -- $0236f
          9072 => x"7b", -- $02370
          9073 => x"7b", -- $02371
          9074 => x"7e", -- $02372
          9075 => x"80", -- $02373
          9076 => x"82", -- $02374
          9077 => x"81", -- $02375
          9078 => x"7f", -- $02376
          9079 => x"7b", -- $02377
          9080 => x"7a", -- $02378
          9081 => x"7a", -- $02379
          9082 => x"7c", -- $0237a
          9083 => x"7e", -- $0237b
          9084 => x"7f", -- $0237c
          9085 => x"7f", -- $0237d
          9086 => x"7f", -- $0237e
          9087 => x"7f", -- $0237f
          9088 => x"80", -- $02380
          9089 => x"81", -- $02381
          9090 => x"82", -- $02382
          9091 => x"84", -- $02383
          9092 => x"84", -- $02384
          9093 => x"83", -- $02385
          9094 => x"83", -- $02386
          9095 => x"84", -- $02387
          9096 => x"86", -- $02388
          9097 => x"87", -- $02389
          9098 => x"88", -- $0238a
          9099 => x"87", -- $0238b
          9100 => x"84", -- $0238c
          9101 => x"83", -- $0238d
          9102 => x"82", -- $0238e
          9103 => x"82", -- $0238f
          9104 => x"82", -- $02390
          9105 => x"82", -- $02391
          9106 => x"83", -- $02392
          9107 => x"83", -- $02393
          9108 => x"85", -- $02394
          9109 => x"86", -- $02395
          9110 => x"86", -- $02396
          9111 => x"82", -- $02397
          9112 => x"81", -- $02398
          9113 => x"7f", -- $02399
          9114 => x"7f", -- $0239a
          9115 => x"81", -- $0239b
          9116 => x"81", -- $0239c
          9117 => x"83", -- $0239d
          9118 => x"82", -- $0239e
          9119 => x"80", -- $0239f
          9120 => x"7f", -- $023a0
          9121 => x"7d", -- $023a1
          9122 => x"7d", -- $023a2
          9123 => x"7e", -- $023a3
          9124 => x"7f", -- $023a4
          9125 => x"7e", -- $023a5
          9126 => x"7d", -- $023a6
          9127 => x"7b", -- $023a7
          9128 => x"7b", -- $023a8
          9129 => x"7d", -- $023a9
          9130 => x"7e", -- $023aa
          9131 => x"80", -- $023ab
          9132 => x"80", -- $023ac
          9133 => x"80", -- $023ad
          9134 => x"7e", -- $023ae
          9135 => x"7e", -- $023af
          9136 => x"7e", -- $023b0
          9137 => x"7f", -- $023b1
          9138 => x"80", -- $023b2
          9139 => x"80", -- $023b3
          9140 => x"81", -- $023b4
          9141 => x"80", -- $023b5
          9142 => x"80", -- $023b6
          9143 => x"7f", -- $023b7
          9144 => x"7f", -- $023b8
          9145 => x"80", -- $023b9
          9146 => x"80", -- $023ba
          9147 => x"81", -- $023bb
          9148 => x"81", -- $023bc
          9149 => x"81", -- $023bd
          9150 => x"82", -- $023be
          9151 => x"82", -- $023bf
          9152 => x"83", -- $023c0
          9153 => x"82", -- $023c1
          9154 => x"82", -- $023c2
          9155 => x"82", -- $023c3
          9156 => x"81", -- $023c4
          9157 => x"81", -- $023c5
          9158 => x"81", -- $023c6
          9159 => x"81", -- $023c7
          9160 => x"81", -- $023c8
          9161 => x"83", -- $023c9
          9162 => x"83", -- $023ca
          9163 => x"83", -- $023cb
          9164 => x"84", -- $023cc
          9165 => x"85", -- $023cd
          9166 => x"86", -- $023ce
          9167 => x"85", -- $023cf
          9168 => x"84", -- $023d0
          9169 => x"83", -- $023d1
          9170 => x"81", -- $023d2
          9171 => x"80", -- $023d3
          9172 => x"80", -- $023d4
          9173 => x"80", -- $023d5
          9174 => x"80", -- $023d6
          9175 => x"82", -- $023d7
          9176 => x"83", -- $023d8
          9177 => x"83", -- $023d9
          9178 => x"83", -- $023da
          9179 => x"83", -- $023db
          9180 => x"83", -- $023dc
          9181 => x"82", -- $023dd
          9182 => x"82", -- $023de
          9183 => x"80", -- $023df
          9184 => x"80", -- $023e0
          9185 => x"80", -- $023e1
          9186 => x"7e", -- $023e2
          9187 => x"80", -- $023e3
          9188 => x"80", -- $023e4
          9189 => x"80", -- $023e5
          9190 => x"80", -- $023e6
          9191 => x"80", -- $023e7
          9192 => x"7f", -- $023e8
          9193 => x"7e", -- $023e9
          9194 => x"7e", -- $023ea
          9195 => x"7f", -- $023eb
          9196 => x"80", -- $023ec
          9197 => x"80", -- $023ed
          9198 => x"80", -- $023ee
          9199 => x"80", -- $023ef
          9200 => x"80", -- $023f0
          9201 => x"80", -- $023f1
          9202 => x"80", -- $023f2
          9203 => x"80", -- $023f3
          9204 => x"80", -- $023f4
          9205 => x"80", -- $023f5
          9206 => x"80", -- $023f6
          9207 => x"80", -- $023f7
          9208 => x"7f", -- $023f8
          9209 => x"80", -- $023f9
          9210 => x"80", -- $023fa
          9211 => x"80", -- $023fb
          9212 => x"80", -- $023fc
          9213 => x"80", -- $023fd
          9214 => x"81", -- $023fe
          9215 => x"81", -- $023ff
          9216 => x"82", -- $02400
          9217 => x"82", -- $02401
          9218 => x"83", -- $02402
          9219 => x"82", -- $02403
          9220 => x"82", -- $02404
          9221 => x"81", -- $02405
          9222 => x"81", -- $02406
          9223 => x"82", -- $02407
          9224 => x"82", -- $02408
          9225 => x"82", -- $02409
          9226 => x"82", -- $0240a
          9227 => x"82", -- $0240b
          9228 => x"81", -- $0240c
          9229 => x"82", -- $0240d
          9230 => x"82", -- $0240e
          9231 => x"83", -- $0240f
          9232 => x"84", -- $02410
          9233 => x"84", -- $02411
          9234 => x"85", -- $02412
          9235 => x"84", -- $02413
          9236 => x"84", -- $02414
          9237 => x"84", -- $02415
          9238 => x"84", -- $02416
          9239 => x"83", -- $02417
          9240 => x"85", -- $02418
          9241 => x"84", -- $02419
          9242 => x"84", -- $0241a
          9243 => x"83", -- $0241b
          9244 => x"82", -- $0241c
          9245 => x"83", -- $0241d
          9246 => x"84", -- $0241e
          9247 => x"84", -- $0241f
          9248 => x"83", -- $02420
          9249 => x"82", -- $02421
          9250 => x"81", -- $02422
          9251 => x"81", -- $02423
          9252 => x"81", -- $02424
          9253 => x"81", -- $02425
          9254 => x"81", -- $02426
          9255 => x"80", -- $02427
          9256 => x"80", -- $02428
          9257 => x"80", -- $02429
          9258 => x"80", -- $0242a
          9259 => x"80", -- $0242b
          9260 => x"80", -- $0242c
          9261 => x"80", -- $0242d
          9262 => x"80", -- $0242e
          9263 => x"80", -- $0242f
          9264 => x"80", -- $02430
          9265 => x"80", -- $02431
          9266 => x"80", -- $02432
          9267 => x"7f", -- $02433
          9268 => x"7e", -- $02434
          9269 => x"7f", -- $02435
          9270 => x"7f", -- $02436
          9271 => x"7f", -- $02437
          9272 => x"7e", -- $02438
          9273 => x"7e", -- $02439
          9274 => x"7e", -- $0243a
          9275 => x"7e", -- $0243b
          9276 => x"7d", -- $0243c
          9277 => x"7e", -- $0243d
          9278 => x"7f", -- $0243e
          9279 => x"7f", -- $0243f
          9280 => x"80", -- $02440
          9281 => x"80", -- $02441
          9282 => x"81", -- $02442
          9283 => x"81", -- $02443
          9284 => x"81", -- $02444
          9285 => x"81", -- $02445
          9286 => x"82", -- $02446
          9287 => x"82", -- $02447
          9288 => x"83", -- $02448
          9289 => x"82", -- $02449
          9290 => x"82", -- $0244a
          9291 => x"82", -- $0244b
          9292 => x"82", -- $0244c
          9293 => x"83", -- $0244d
          9294 => x"83", -- $0244e
          9295 => x"83", -- $0244f
          9296 => x"82", -- $02450
          9297 => x"83", -- $02451
          9298 => x"83", -- $02452
          9299 => x"82", -- $02453
          9300 => x"82", -- $02454
          9301 => x"82", -- $02455
          9302 => x"83", -- $02456
          9303 => x"83", -- $02457
          9304 => x"82", -- $02458
          9305 => x"82", -- $02459
          9306 => x"82", -- $0245a
          9307 => x"81", -- $0245b
          9308 => x"81", -- $0245c
          9309 => x"80", -- $0245d
          9310 => x"80", -- $0245e
          9311 => x"80", -- $0245f
          9312 => x"80", -- $02460
          9313 => x"80", -- $02461
          9314 => x"80", -- $02462
          9315 => x"7f", -- $02463
          9316 => x"7f", -- $02464
          9317 => x"7e", -- $02465
          9318 => x"7e", -- $02466
          9319 => x"7f", -- $02467
          9320 => x"7f", -- $02468
          9321 => x"7f", -- $02469
          9322 => x"7f", -- $0246a
          9323 => x"7f", -- $0246b
          9324 => x"7e", -- $0246c
          9325 => x"7e", -- $0246d
          9326 => x"7e", -- $0246e
          9327 => x"7e", -- $0246f
          9328 => x"7e", -- $02470
          9329 => x"7e", -- $02471
          9330 => x"7e", -- $02472
          9331 => x"7d", -- $02473
          9332 => x"7d", -- $02474
          9333 => x"7d", -- $02475
          9334 => x"7d", -- $02476
          9335 => x"7d", -- $02477
          9336 => x"7d", -- $02478
          9337 => x"7d", -- $02479
          9338 => x"7d", -- $0247a
          9339 => x"7e", -- $0247b
          9340 => x"7e", -- $0247c
          9341 => x"7e", -- $0247d
          9342 => x"7f", -- $0247e
          9343 => x"7f", -- $0247f
          9344 => x"80", -- $02480
          9345 => x"80", -- $02481
          9346 => x"80", -- $02482
          9347 => x"80", -- $02483
          9348 => x"80", -- $02484
          9349 => x"80", -- $02485
          9350 => x"80", -- $02486
          9351 => x"80", -- $02487
          9352 => x"80", -- $02488
          9353 => x"80", -- $02489
          9354 => x"80", -- $0248a
          9355 => x"80", -- $0248b
          9356 => x"80", -- $0248c
          9357 => x"81", -- $0248d
          9358 => x"81", -- $0248e
          9359 => x"81", -- $0248f
          9360 => x"82", -- $02490
          9361 => x"81", -- $02491
          9362 => x"81", -- $02492
          9363 => x"81", -- $02493
          9364 => x"81", -- $02494
          9365 => x"81", -- $02495
          9366 => x"81", -- $02496
          9367 => x"81", -- $02497
          9368 => x"81", -- $02498
          9369 => x"81", -- $02499
          9370 => x"80", -- $0249a
          9371 => x"80", -- $0249b
          9372 => x"80", -- $0249c
          9373 => x"80", -- $0249d
          9374 => x"80", -- $0249e
          9375 => x"80", -- $0249f
          9376 => x"7f", -- $024a0
          9377 => x"7f", -- $024a1
          9378 => x"7e", -- $024a2
          9379 => x"7e", -- $024a3
          9380 => x"7f", -- $024a4
          9381 => x"7f", -- $024a5
          9382 => x"7f", -- $024a6
          9383 => x"7f", -- $024a7
          9384 => x"7e", -- $024a8
          9385 => x"7e", -- $024a9
          9386 => x"7e", -- $024aa
          9387 => x"7d", -- $024ab
          9388 => x"7d", -- $024ac
          9389 => x"7d", -- $024ad
          9390 => x"7d", -- $024ae
          9391 => x"7d", -- $024af
          9392 => x"7e", -- $024b0
          9393 => x"7e", -- $024b1
          9394 => x"7e", -- $024b2
          9395 => x"7e", -- $024b3
          9396 => x"7e", -- $024b4
          9397 => x"7e", -- $024b5
          9398 => x"7e", -- $024b6
          9399 => x"7e", -- $024b7
          9400 => x"7f", -- $024b8
          9401 => x"7f", -- $024b9
          9402 => x"7f", -- $024ba
          9403 => x"80", -- $024bb
          9404 => x"80", -- $024bc
          9405 => x"80", -- $024bd
          9406 => x"80", -- $024be
          9407 => x"80", -- $024bf
          9408 => x"80", -- $024c0
          9409 => x"80", -- $024c1
          9410 => x"80", -- $024c2
          9411 => x"80", -- $024c3
          9412 => x"80", -- $024c4
          9413 => x"81", -- $024c5
          9414 => x"81", -- $024c6
          9415 => x"81", -- $024c7
          9416 => x"81", -- $024c8
          9417 => x"81", -- $024c9
          9418 => x"81", -- $024ca
          9419 => x"80", -- $024cb
          9420 => x"81", -- $024cc
          9421 => x"81", -- $024cd
          9422 => x"81", -- $024ce
          9423 => x"81", -- $024cf
          9424 => x"81", -- $024d0
          9425 => x"81", -- $024d1
          9426 => x"80", -- $024d2
          9427 => x"80", -- $024d3
          9428 => x"80", -- $024d4
          9429 => x"80", -- $024d5
          9430 => x"80", -- $024d6
          9431 => x"80", -- $024d7
          9432 => x"80", -- $024d8
          9433 => x"80", -- $024d9
          9434 => x"80", -- $024da
          9435 => x"80", -- $024db
          9436 => x"7f", -- $024dc
          9437 => x"7f", -- $024dd
          9438 => x"7f", -- $024de
          9439 => x"7f", -- $024df
          9440 => x"7f", -- $024e0
          9441 => x"7f", -- $024e1
          9442 => x"7f", -- $024e2
          9443 => x"7e", -- $024e3
          9444 => x"7f", -- $024e4
          9445 => x"7e", -- $024e5
          9446 => x"7e", -- $024e6
          9447 => x"7e", -- $024e7
          9448 => x"7e", -- $024e8
          9449 => x"7e", -- $024e9
          9450 => x"7e", -- $024ea
          9451 => x"7e", -- $024eb
          9452 => x"7e", -- $024ec
          9453 => x"7e", -- $024ed
          9454 => x"7e", -- $024ee
          9455 => x"7e", -- $024ef
          9456 => x"7e", -- $024f0
          9457 => x"7e", -- $024f1
          9458 => x"7e", -- $024f2
          9459 => x"7e", -- $024f3
          9460 => x"7f", -- $024f4
          9461 => x"7f", -- $024f5
          9462 => x"7f", -- $024f6
          9463 => x"7f", -- $024f7
          9464 => x"7f", -- $024f8
          9465 => x"7f", -- $024f9
          9466 => x"7f", -- $024fa
          9467 => x"7f", -- $024fb
          9468 => x"80", -- $024fc
          9469 => x"80", -- $024fd
          9470 => x"80", -- $024fe
          9471 => x"80", -- $024ff
          9472 => x"80", -- $02500
          9473 => x"80", -- $02501
          9474 => x"80", -- $02502
          9475 => x"80", -- $02503
          9476 => x"80", -- $02504
          9477 => x"80", -- $02505
          9478 => x"80", -- $02506
          9479 => x"80", -- $02507
          9480 => x"80", -- $02508
          9481 => x"80", -- $02509
          9482 => x"80", -- $0250a
          9483 => x"80", -- $0250b
          9484 => x"80", -- $0250c
          9485 => x"7f", -- $0250d
          9486 => x"80", -- $0250e
          9487 => x"80", -- $0250f
          9488 => x"80", -- $02510
          9489 => x"80", -- $02511
          9490 => x"80", -- $02512
          9491 => x"80", -- $02513
          9492 => x"80", -- $02514
          9493 => x"80", -- $02515
          9494 => x"80", -- $02516
          9495 => x"80", -- $02517
          9496 => x"80", -- $02518
          9497 => x"80", -- $02519
          9498 => x"80", -- $0251a
          9499 => x"80", -- $0251b
          9500 => x"80", -- $0251c
          9501 => x"7f", -- $0251d
          9502 => x"7f", -- $0251e
          9503 => x"7f", -- $0251f
          9504 => x"7e", -- $02520
          9505 => x"7e", -- $02521
          9506 => x"7e", -- $02522
          9507 => x"7e", -- $02523
          9508 => x"7e", -- $02524
          9509 => x"7d", -- $02525
          9510 => x"7d", -- $02526
          9511 => x"7d", -- $02527
          9512 => x"7d", -- $02528
          9513 => x"7c", -- $02529
          9514 => x"7d", -- $0252a
          9515 => x"7e", -- $0252b
          9516 => x"7e", -- $0252c
          9517 => x"7e", -- $0252d
          9518 => x"7e", -- $0252e
          9519 => x"7e", -- $0252f
          9520 => x"7e", -- $02530
          9521 => x"7e", -- $02531
          9522 => x"7e", -- $02532
          9523 => x"7e", -- $02533
          9524 => x"7e", -- $02534
          9525 => x"7e", -- $02535
          9526 => x"7e", -- $02536
          9527 => x"7f", -- $02537
          9528 => x"7f", -- $02538
          9529 => x"7f", -- $02539
          9530 => x"7f", -- $0253a
          9531 => x"80", -- $0253b
          9532 => x"7f", -- $0253c
          9533 => x"7f", -- $0253d
          9534 => x"7f", -- $0253e
          9535 => x"7e", -- $0253f
          9536 => x"7e", -- $02540
          9537 => x"7d", -- $02541
          9538 => x"7e", -- $02542
          9539 => x"7f", -- $02543
          9540 => x"80", -- $02544
          9541 => x"7f", -- $02545
          9542 => x"7f", -- $02546
          9543 => x"7f", -- $02547
          9544 => x"80", -- $02548
          9545 => x"80", -- $02549
          9546 => x"80", -- $0254a
          9547 => x"80", -- $0254b
          9548 => x"80", -- $0254c
          9549 => x"80", -- $0254d
          9550 => x"80", -- $0254e
          9551 => x"80", -- $0254f
          9552 => x"80", -- $02550
          9553 => x"80", -- $02551
          9554 => x"80", -- $02552
          9555 => x"80", -- $02553
          9556 => x"80", -- $02554
          9557 => x"80", -- $02555
          9558 => x"80", -- $02556
          9559 => x"7f", -- $02557
          9560 => x"7f", -- $02558
          9561 => x"7f", -- $02559
          9562 => x"7f", -- $0255a
          9563 => x"7f", -- $0255b
          9564 => x"7f", -- $0255c
          9565 => x"7f", -- $0255d
          9566 => x"7f", -- $0255e
          9567 => x"7f", -- $0255f
          9568 => x"7f", -- $02560
          9569 => x"7e", -- $02561
          9570 => x"7e", -- $02562
          9571 => x"7d", -- $02563
          9572 => x"7d", -- $02564
          9573 => x"7e", -- $02565
          9574 => x"7f", -- $02566
          9575 => x"7f", -- $02567
          9576 => x"7f", -- $02568
          9577 => x"7f", -- $02569
          9578 => x"7f", -- $0256a
          9579 => x"7e", -- $0256b
          9580 => x"7e", -- $0256c
          9581 => x"7f", -- $0256d
          9582 => x"7f", -- $0256e
          9583 => x"7f", -- $0256f
          9584 => x"7e", -- $02570
          9585 => x"7f", -- $02571
          9586 => x"7f", -- $02572
          9587 => x"7f", -- $02573
          9588 => x"80", -- $02574
          9589 => x"80", -- $02575
          9590 => x"80", -- $02576
          9591 => x"80", -- $02577
          9592 => x"80", -- $02578
          9593 => x"7f", -- $02579
          9594 => x"7f", -- $0257a
          9595 => x"80", -- $0257b
          9596 => x"80", -- $0257c
          9597 => x"80", -- $0257d
          9598 => x"80", -- $0257e
          9599 => x"80", -- $0257f
          9600 => x"80", -- $02580
          9601 => x"80", -- $02581
          9602 => x"80", -- $02582
          9603 => x"80", -- $02583
          9604 => x"80", -- $02584
          9605 => x"80", -- $02585
          9606 => x"80", -- $02586
          9607 => x"80", -- $02587
          9608 => x"80", -- $02588
          9609 => x"7f", -- $02589
          9610 => x"80", -- $0258a
          9611 => x"80", -- $0258b
          9612 => x"80", -- $0258c
          9613 => x"80", -- $0258d
          9614 => x"80", -- $0258e
          9615 => x"80", -- $0258f
          9616 => x"80", -- $02590
          9617 => x"7f", -- $02591
          9618 => x"7f", -- $02592
          9619 => x"7f", -- $02593
          9620 => x"7f", -- $02594
          9621 => x"80", -- $02595
          9622 => x"80", -- $02596
          9623 => x"80", -- $02597
          9624 => x"7f", -- $02598
          9625 => x"80", -- $02599
          9626 => x"7f", -- $0259a
          9627 => x"7f", -- $0259b
          9628 => x"7f", -- $0259c
          9629 => x"7f", -- $0259d
          9630 => x"7f", -- $0259e
          9631 => x"7e", -- $0259f
          9632 => x"7f", -- $025a0
          9633 => x"7e", -- $025a1
          9634 => x"7e", -- $025a2
          9635 => x"7f", -- $025a3
          9636 => x"7e", -- $025a4
          9637 => x"80", -- $025a5
          9638 => x"7f", -- $025a6
          9639 => x"7f", -- $025a7
          9640 => x"7f", -- $025a8
          9641 => x"80", -- $025a9
          9642 => x"7f", -- $025aa
          9643 => x"80", -- $025ab
          9644 => x"80", -- $025ac
          9645 => x"80", -- $025ad
          9646 => x"80", -- $025ae
          9647 => x"80", -- $025af
          9648 => x"81", -- $025b0
          9649 => x"7f", -- $025b1
          9650 => x"7f", -- $025b2
          9651 => x"7e", -- $025b3
          9652 => x"80", -- $025b4
          9653 => x"81", -- $025b5
          9654 => x"81", -- $025b6
          9655 => x"80", -- $025b7
          9656 => x"80", -- $025b8
          9657 => x"7f", -- $025b9
          9658 => x"80", -- $025ba
          9659 => x"80", -- $025bb
          9660 => x"7f", -- $025bc
          9661 => x"80", -- $025bd
          9662 => x"80", -- $025be
          9663 => x"81", -- $025bf
          9664 => x"80", -- $025c0
          9665 => x"81", -- $025c1
          9666 => x"7f", -- $025c2
          9667 => x"82", -- $025c3
          9668 => x"80", -- $025c4
          9669 => x"82", -- $025c5
          9670 => x"80", -- $025c6
          9671 => x"80", -- $025c7
          9672 => x"80", -- $025c8
          9673 => x"80", -- $025c9
          9674 => x"80", -- $025ca
          9675 => x"80", -- $025cb
          9676 => x"81", -- $025cc
          9677 => x"7f", -- $025cd
          9678 => x"81", -- $025ce
          9679 => x"7e", -- $025cf
          9680 => x"80", -- $025d0
          9681 => x"7f", -- $025d1
          9682 => x"80", -- $025d2
          9683 => x"80", -- $025d3
          9684 => x"80", -- $025d4
          9685 => x"7f", -- $025d5
          9686 => x"80", -- $025d6
          9687 => x"80", -- $025d7
          9688 => x"80", -- $025d8
          9689 => x"80", -- $025d9
          9690 => x"80", -- $025da
          9691 => x"80", -- $025db
          9692 => x"7f", -- $025dc
          9693 => x"80", -- $025dd
          9694 => x"7f", -- $025de
          9695 => x"80", -- $025df
          9696 => x"7e", -- $025e0
          9697 => x"80", -- $025e1
          9698 => x"7e", -- $025e2
          9699 => x"80", -- $025e3
          9700 => x"7e", -- $025e4
          9701 => x"80", -- $025e5
          9702 => x"7e", -- $025e6
          9703 => x"80", -- $025e7
          9704 => x"7f", -- $025e8
          9705 => x"80", -- $025e9
          9706 => x"80", -- $025ea
          9707 => x"80", -- $025eb
          9708 => x"80", -- $025ec
          9709 => x"80", -- $025ed
          9710 => x"82", -- $025ee
          9711 => x"7f", -- $025ef
          9712 => x"82", -- $025f0
          9713 => x"7e", -- $025f1
          9714 => x"81", -- $025f2
          9715 => x"80", -- $025f3
          9716 => x"80", -- $025f4
          9717 => x"80", -- $025f5
          9718 => x"80", -- $025f6
          9719 => x"80", -- $025f7
          9720 => x"80", -- $025f8
          9721 => x"80", -- $025f9
          9722 => x"7f", -- $025fa
          9723 => x"80", -- $025fb
          9724 => x"80", -- $025fc
          9725 => x"80", -- $025fd
          9726 => x"81", -- $025fe
          9727 => x"81", -- $025ff
          9728 => x"80", -- $02600
          9729 => x"82", -- $02601
          9730 => x"80", -- $02602
          9731 => x"82", -- $02603
          9732 => x"81", -- $02604
          9733 => x"81", -- $02605
          9734 => x"81", -- $02606
          9735 => x"81", -- $02607
          9736 => x"81", -- $02608
          9737 => x"82", -- $02609
          9738 => x"80", -- $0260a
          9739 => x"81", -- $0260b
          9740 => x"81", -- $0260c
          9741 => x"80", -- $0260d
          9742 => x"80", -- $0260e
          9743 => x"80", -- $0260f
          9744 => x"81", -- $02610
          9745 => x"80", -- $02611
          9746 => x"81", -- $02612
          9747 => x"80", -- $02613
          9748 => x"82", -- $02614
          9749 => x"80", -- $02615
          9750 => x"82", -- $02616
          9751 => x"82", -- $02617
          9752 => x"7f", -- $02618
          9753 => x"81", -- $02619
          9754 => x"80", -- $0261a
          9755 => x"80", -- $0261b
          9756 => x"80", -- $0261c
          9757 => x"80", -- $0261d
          9758 => x"7f", -- $0261e
          9759 => x"81", -- $0261f
          9760 => x"7f", -- $02620
          9761 => x"80", -- $02621
          9762 => x"80", -- $02622
          9763 => x"7f", -- $02623
          9764 => x"80", -- $02624
          9765 => x"80", -- $02625
          9766 => x"80", -- $02626
          9767 => x"80", -- $02627
          9768 => x"80", -- $02628
          9769 => x"7f", -- $02629
          9770 => x"81", -- $0262a
          9771 => x"7f", -- $0262b
          9772 => x"81", -- $0262c
          9773 => x"80", -- $0262d
          9774 => x"80", -- $0262e
          9775 => x"81", -- $0262f
          9776 => x"80", -- $02630
          9777 => x"80", -- $02631
          9778 => x"7f", -- $02632
          9779 => x"80", -- $02633
          9780 => x"80", -- $02634
          9781 => x"81", -- $02635
          9782 => x"7f", -- $02636
          9783 => x"82", -- $02637
          9784 => x"80", -- $02638
          9785 => x"81", -- $02639
          9786 => x"82", -- $0263a
          9787 => x"80", -- $0263b
          9788 => x"82", -- $0263c
          9789 => x"80", -- $0263d
          9790 => x"81", -- $0263e
          9791 => x"82", -- $0263f
          9792 => x"80", -- $02640
          9793 => x"82", -- $02641
          9794 => x"80", -- $02642
          9795 => x"81", -- $02643
          9796 => x"80", -- $02644
          9797 => x"81", -- $02645
          9798 => x"80", -- $02646
          9799 => x"81", -- $02647
          9800 => x"81", -- $02648
          9801 => x"7e", -- $02649
          9802 => x"82", -- $0264a
          9803 => x"80", -- $0264b
          9804 => x"81", -- $0264c
          9805 => x"80", -- $0264d
          9806 => x"7f", -- $0264e
          9807 => x"80", -- $0264f
          9808 => x"80", -- $02650
          9809 => x"80", -- $02651
          9810 => x"81", -- $02652
          9811 => x"81", -- $02653
          9812 => x"80", -- $02654
          9813 => x"83", -- $02655
          9814 => x"80", -- $02656
          9815 => x"81", -- $02657
          9816 => x"80", -- $02658
          9817 => x"80", -- $02659
          9818 => x"80", -- $0265a
          9819 => x"80", -- $0265b
          9820 => x"80", -- $0265c
          9821 => x"80", -- $0265d
          9822 => x"80", -- $0265e
          9823 => x"80", -- $0265f
          9824 => x"82", -- $02660
          9825 => x"80", -- $02661
          9826 => x"82", -- $02662
          9827 => x"81", -- $02663
          9828 => x"81", -- $02664
          9829 => x"83", -- $02665
          9830 => x"81", -- $02666
          9831 => x"81", -- $02667
          9832 => x"81", -- $02668
          9833 => x"81", -- $02669
          9834 => x"81", -- $0266a
          9835 => x"83", -- $0266b
          9836 => x"80", -- $0266c
          9837 => x"81", -- $0266d
          9838 => x"81", -- $0266e
          9839 => x"80", -- $0266f
          9840 => x"82", -- $02670
          9841 => x"81", -- $02671
          9842 => x"80", -- $02672
          9843 => x"80", -- $02673
          9844 => x"81", -- $02674
          9845 => x"81", -- $02675
          9846 => x"84", -- $02676
          9847 => x"82", -- $02677
          9848 => x"82", -- $02678
          9849 => x"82", -- $02679
          9850 => x"80", -- $0267a
          9851 => x"83", -- $0267b
          9852 => x"81", -- $0267c
          9853 => x"80", -- $0267d
          9854 => x"81", -- $0267e
          9855 => x"80", -- $0267f
          9856 => x"82", -- $02680
          9857 => x"82", -- $02681
          9858 => x"81", -- $02682
          9859 => x"81", -- $02683
          9860 => x"81", -- $02684
          9861 => x"81", -- $02685
          9862 => x"82", -- $02686
          9863 => x"83", -- $02687
          9864 => x"81", -- $02688
          9865 => x"81", -- $02689
          9866 => x"80", -- $0268a
          9867 => x"80", -- $0268b
          9868 => x"82", -- $0268c
          9869 => x"80", -- $0268d
          9870 => x"80", -- $0268e
          9871 => x"81", -- $0268f
          9872 => x"81", -- $02690
          9873 => x"82", -- $02691
          9874 => x"82", -- $02692
          9875 => x"81", -- $02693
          9876 => x"80", -- $02694
          9877 => x"82", -- $02695
          9878 => x"81", -- $02696
          9879 => x"82", -- $02697
          9880 => x"81", -- $02698
          9881 => x"81", -- $02699
          9882 => x"81", -- $0269a
          9883 => x"81", -- $0269b
          9884 => x"81", -- $0269c
          9885 => x"81", -- $0269d
          9886 => x"81", -- $0269e
          9887 => x"80", -- $0269f
          9888 => x"81", -- $026a0
          9889 => x"80", -- $026a1
          9890 => x"80", -- $026a2
          9891 => x"80", -- $026a3
          9892 => x"80", -- $026a4
          9893 => x"81", -- $026a5
          9894 => x"82", -- $026a6
          9895 => x"81", -- $026a7
          9896 => x"82", -- $026a8
          9897 => x"82", -- $026a9
          9898 => x"82", -- $026aa
          9899 => x"83", -- $026ab
          9900 => x"83", -- $026ac
          9901 => x"83", -- $026ad
          9902 => x"82", -- $026ae
          9903 => x"82", -- $026af
          9904 => x"82", -- $026b0
          9905 => x"82", -- $026b1
          9906 => x"82", -- $026b2
          9907 => x"81", -- $026b3
          9908 => x"80", -- $026b4
          9909 => x"82", -- $026b5
          9910 => x"82", -- $026b6
          9911 => x"83", -- $026b7
          9912 => x"82", -- $026b8
          9913 => x"81", -- $026b9
          9914 => x"82", -- $026ba
          9915 => x"81", -- $026bb
          9916 => x"82", -- $026bc
          9917 => x"81", -- $026bd
          9918 => x"81", -- $026be
          9919 => x"81", -- $026bf
          9920 => x"84", -- $026c0
          9921 => x"84", -- $026c1
          9922 => x"82", -- $026c2
          9923 => x"82", -- $026c3
          9924 => x"81", -- $026c4
          9925 => x"82", -- $026c5
          9926 => x"82", -- $026c6
          9927 => x"82", -- $026c7
          9928 => x"81", -- $026c8
          9929 => x"80", -- $026c9
          9930 => x"81", -- $026ca
          9931 => x"82", -- $026cb
          9932 => x"82", -- $026cc
          9933 => x"82", -- $026cd
          9934 => x"81", -- $026ce
          9935 => x"81", -- $026cf
          9936 => x"81", -- $026d0
          9937 => x"82", -- $026d1
          9938 => x"80", -- $026d2
          9939 => x"80", -- $026d3
          9940 => x"80", -- $026d4
          9941 => x"80", -- $026d5
          9942 => x"82", -- $026d6
          9943 => x"81", -- $026d7
          9944 => x"80", -- $026d8
          9945 => x"80", -- $026d9
          9946 => x"80", -- $026da
          9947 => x"81", -- $026db
          9948 => x"81", -- $026dc
          9949 => x"80", -- $026dd
          9950 => x"7f", -- $026de
          9951 => x"80", -- $026df
          9952 => x"80", -- $026e0
          9953 => x"80", -- $026e1
          9954 => x"80", -- $026e2
          9955 => x"80", -- $026e3
          9956 => x"80", -- $026e4
          9957 => x"81", -- $026e5
          9958 => x"81", -- $026e6
          9959 => x"81", -- $026e7
          9960 => x"80", -- $026e8
          9961 => x"80", -- $026e9
          9962 => x"80", -- $026ea
          9963 => x"81", -- $026eb
          9964 => x"80", -- $026ec
          9965 => x"80", -- $026ed
          9966 => x"81", -- $026ee
          9967 => x"81", -- $026ef
          9968 => x"83", -- $026f0
          9969 => x"82", -- $026f1
          9970 => x"82", -- $026f2
          9971 => x"82", -- $026f3
          9972 => x"81", -- $026f4
          9973 => x"82", -- $026f5
          9974 => x"82", -- $026f6
          9975 => x"82", -- $026f7
          9976 => x"82", -- $026f8
          9977 => x"83", -- $026f9
          9978 => x"83", -- $026fa
          9979 => x"83", -- $026fb
          9980 => x"83", -- $026fc
          9981 => x"82", -- $026fd
          9982 => x"82", -- $026fe
          9983 => x"82", -- $026ff
          9984 => x"83", -- $02700
          9985 => x"84", -- $02701
          9986 => x"83", -- $02702
          9987 => x"83", -- $02703
          9988 => x"82", -- $02704
          9989 => x"82", -- $02705
          9990 => x"82", -- $02706
          9991 => x"81", -- $02707
          9992 => x"80", -- $02708
          9993 => x"80", -- $02709
          9994 => x"7f", -- $0270a
          9995 => x"7f", -- $0270b
          9996 => x"7e", -- $0270c
          9997 => x"7d", -- $0270d
          9998 => x"7c", -- $0270e
          9999 => x"7c", -- $0270f
          10000 => x"7b", -- $02710
          10001 => x"7a", -- $02711
          10002 => x"7a", -- $02712
          10003 => x"7b", -- $02713
          10004 => x"7b", -- $02714
          10005 => x"7c", -- $02715
          10006 => x"7e", -- $02716
          10007 => x"7f", -- $02717
          10008 => x"80", -- $02718
          10009 => x"80", -- $02719
          10010 => x"80", -- $0271a
          10011 => x"80", -- $0271b
          10012 => x"80", -- $0271c
          10013 => x"81", -- $0271d
          10014 => x"80", -- $0271e
          10015 => x"81", -- $0271f
          10016 => x"82", -- $02720
          10017 => x"82", -- $02721
          10018 => x"82", -- $02722
          10019 => x"84", -- $02723
          10020 => x"85", -- $02724
          10021 => x"85", -- $02725
          10022 => x"86", -- $02726
          10023 => x"86", -- $02727
          10024 => x"86", -- $02728
          10025 => x"87", -- $02729
          10026 => x"86", -- $0272a
          10027 => x"86", -- $0272b
          10028 => x"85", -- $0272c
          10029 => x"83", -- $0272d
          10030 => x"83", -- $0272e
          10031 => x"83", -- $0272f
          10032 => x"82", -- $02730
          10033 => x"81", -- $02731
          10034 => x"81", -- $02732
          10035 => x"80", -- $02733
          10036 => x"81", -- $02734
          10037 => x"80", -- $02735
          10038 => x"80", -- $02736
          10039 => x"80", -- $02737
          10040 => x"7f", -- $02738
          10041 => x"7f", -- $02739
          10042 => x"7f", -- $0273a
          10043 => x"7e", -- $0273b
          10044 => x"7d", -- $0273c
          10045 => x"7d", -- $0273d
          10046 => x"7d", -- $0273e
          10047 => x"7d", -- $0273f
          10048 => x"7e", -- $02740
          10049 => x"7f", -- $02741
          10050 => x"7f", -- $02742
          10051 => x"80", -- $02743
          10052 => x"81", -- $02744
          10053 => x"83", -- $02745
          10054 => x"84", -- $02746
          10055 => x"84", -- $02747
          10056 => x"84", -- $02748
          10057 => x"84", -- $02749
          10058 => x"83", -- $0274a
          10059 => x"82", -- $0274b
          10060 => x"81", -- $0274c
          10061 => x"80", -- $0274d
          10062 => x"7e", -- $0274e
          10063 => x"7c", -- $0274f
          10064 => x"7b", -- $02750
          10065 => x"78", -- $02751
          10066 => x"79", -- $02752
          10067 => x"7a", -- $02753
          10068 => x"7b", -- $02754
          10069 => x"7d", -- $02755
          10070 => x"7e", -- $02756
          10071 => x"7f", -- $02757
          10072 => x"80", -- $02758
          10073 => x"80", -- $02759
          10074 => x"80", -- $0275a
          10075 => x"7f", -- $0275b
          10076 => x"7f", -- $0275c
          10077 => x"7d", -- $0275d
          10078 => x"7e", -- $0275e
          10079 => x"7e", -- $0275f
          10080 => x"7e", -- $02760
          10081 => x"7e", -- $02761
          10082 => x"7e", -- $02762
          10083 => x"80", -- $02763
          10084 => x"80", -- $02764
          10085 => x"81", -- $02765
          10086 => x"83", -- $02766
          10087 => x"84", -- $02767
          10088 => x"85", -- $02768
          10089 => x"86", -- $02769
          10090 => x"87", -- $0276a
          10091 => x"87", -- $0276b
          10092 => x"86", -- $0276c
          10093 => x"85", -- $0276d
          10094 => x"85", -- $0276e
          10095 => x"84", -- $0276f
          10096 => x"83", -- $02770
          10097 => x"83", -- $02771
          10098 => x"82", -- $02772
          10099 => x"82", -- $02773
          10100 => x"82", -- $02774
          10101 => x"81", -- $02775
          10102 => x"80", -- $02776
          10103 => x"81", -- $02777
          10104 => x"81", -- $02778
          10105 => x"82", -- $02779
          10106 => x"82", -- $0277a
          10107 => x"82", -- $0277b
          10108 => x"81", -- $0277c
          10109 => x"80", -- $0277d
          10110 => x"80", -- $0277e
          10111 => x"7f", -- $0277f
          10112 => x"7e", -- $02780
          10113 => x"7c", -- $02781
          10114 => x"7b", -- $02782
          10115 => x"7b", -- $02783
          10116 => x"7b", -- $02784
          10117 => x"7c", -- $02785
          10118 => x"7d", -- $02786
          10119 => x"7e", -- $02787
          10120 => x"7f", -- $02788
          10121 => x"80", -- $02789
          10122 => x"80", -- $0278a
          10123 => x"81", -- $0278b
          10124 => x"81", -- $0278c
          10125 => x"80", -- $0278d
          10126 => x"80", -- $0278e
          10127 => x"80", -- $0278f
          10128 => x"7e", -- $02790
          10129 => x"7d", -- $02791
          10130 => x"7b", -- $02792
          10131 => x"79", -- $02793
          10132 => x"77", -- $02794
          10133 => x"77", -- $02795
          10134 => x"78", -- $02796
          10135 => x"7a", -- $02797
          10136 => x"7c", -- $02798
          10137 => x"7d", -- $02799
          10138 => x"7d", -- $0279a
          10139 => x"7e", -- $0279b
          10140 => x"80", -- $0279c
          10141 => x"80", -- $0279d
          10142 => x"80", -- $0279e
          10143 => x"7f", -- $0279f
          10144 => x"7e", -- $027a0
          10145 => x"7e", -- $027a1
          10146 => x"7f", -- $027a2
          10147 => x"7f", -- $027a3
          10148 => x"7f", -- $027a4
          10149 => x"7f", -- $027a5
          10150 => x"80", -- $027a6
          10151 => x"81", -- $027a7
          10152 => x"84", -- $027a8
          10153 => x"85", -- $027a9
          10154 => x"87", -- $027aa
          10155 => x"89", -- $027ab
          10156 => x"88", -- $027ac
          10157 => x"86", -- $027ad
          10158 => x"84", -- $027ae
          10159 => x"81", -- $027af
          10160 => x"81", -- $027b0
          10161 => x"83", -- $027b1
          10162 => x"81", -- $027b2
          10163 => x"81", -- $027b3
          10164 => x"80", -- $027b4
          10165 => x"80", -- $027b5
          10166 => x"80", -- $027b6
          10167 => x"80", -- $027b7
          10168 => x"80", -- $027b8
          10169 => x"7d", -- $027b9
          10170 => x"7c", -- $027ba
          10171 => x"7b", -- $027bb
          10172 => x"7c", -- $027bc
          10173 => x"7c", -- $027bd
          10174 => x"7c", -- $027be
          10175 => x"7c", -- $027bf
          10176 => x"7d", -- $027c0
          10177 => x"7f", -- $027c1
          10178 => x"81", -- $027c2
          10179 => x"82", -- $027c3
          10180 => x"81", -- $027c4
          10181 => x"81", -- $027c5
          10182 => x"83", -- $027c6
          10183 => x"84", -- $027c7
          10184 => x"84", -- $027c8
          10185 => x"83", -- $027c9
          10186 => x"80", -- $027ca
          10187 => x"7f", -- $027cb
          10188 => x"7d", -- $027cc
          10189 => x"7c", -- $027cd
          10190 => x"7a", -- $027ce
          10191 => x"79", -- $027cf
          10192 => x"77", -- $027d0
          10193 => x"77", -- $027d1
          10194 => x"78", -- $027d2
          10195 => x"79", -- $027d3
          10196 => x"7b", -- $027d4
          10197 => x"7c", -- $027d5
          10198 => x"7d", -- $027d6
          10199 => x"7f", -- $027d7
          10200 => x"80", -- $027d8
          10201 => x"81", -- $027d9
          10202 => x"80", -- $027da
          10203 => x"7f", -- $027db
          10204 => x"7d", -- $027dc
          10205 => x"7c", -- $027dd
          10206 => x"7b", -- $027de
          10207 => x"7a", -- $027df
          10208 => x"79", -- $027e0
          10209 => x"79", -- $027e1
          10210 => x"79", -- $027e2
          10211 => x"7b", -- $027e3
          10212 => x"7d", -- $027e4
          10213 => x"80", -- $027e5
          10214 => x"81", -- $027e6
          10215 => x"83", -- $027e7
          10216 => x"84", -- $027e8
          10217 => x"85", -- $027e9
          10218 => x"85", -- $027ea
          10219 => x"85", -- $027eb
          10220 => x"84", -- $027ec
          10221 => x"82", -- $027ed
          10222 => x"80", -- $027ee
          10223 => x"80", -- $027ef
          10224 => x"7f", -- $027f0
          10225 => x"7e", -- $027f1
          10226 => x"7e", -- $027f2
          10227 => x"7e", -- $027f3
          10228 => x"7f", -- $027f4
          10229 => x"80", -- $027f5
          10230 => x"81", -- $027f6
          10231 => x"82", -- $027f7
          10232 => x"83", -- $027f8
          10233 => x"83", -- $027f9
          10234 => x"84", -- $027fa
          10235 => x"83", -- $027fb
          10236 => x"82", -- $027fc
          10237 => x"82", -- $027fd
          10238 => x"80", -- $027fe
          10239 => x"7f", -- $027ff
          10240 => x"7e", -- $02800
          10241 => x"7d", -- $02801
          10242 => x"7d", -- $02802
          10243 => x"7d", -- $02803
          10244 => x"7c", -- $02804
          10245 => x"7d", -- $02805
          10246 => x"7e", -- $02806
          10247 => x"7f", -- $02807
          10248 => x"80", -- $02808
          10249 => x"80", -- $02809
          10250 => x"80", -- $0280a
          10251 => x"80", -- $0280b
          10252 => x"80", -- $0280c
          10253 => x"7f", -- $0280d
          10254 => x"7e", -- $0280e
          10255 => x"7d", -- $0280f
          10256 => x"7b", -- $02810
          10257 => x"7a", -- $02811
          10258 => x"7a", -- $02812
          10259 => x"7a", -- $02813
          10260 => x"7a", -- $02814
          10261 => x"7b", -- $02815
          10262 => x"7c", -- $02816
          10263 => x"7e", -- $02817
          10264 => x"80", -- $02818
          10265 => x"80", -- $02819
          10266 => x"81", -- $0281a
          10267 => x"81", -- $0281b
          10268 => x"81", -- $0281c
          10269 => x"80", -- $0281d
          10270 => x"80", -- $0281e
          10271 => x"7f", -- $0281f
          10272 => x"7e", -- $02820
          10273 => x"7c", -- $02821
          10274 => x"7c", -- $02822
          10275 => x"7b", -- $02823
          10276 => x"7b", -- $02824
          10277 => x"7b", -- $02825
          10278 => x"7d", -- $02826
          10279 => x"7f", -- $02827
          10280 => x"80", -- $02828
          10281 => x"82", -- $02829
          10282 => x"83", -- $0282a
          10283 => x"84", -- $0282b
          10284 => x"85", -- $0282c
          10285 => x"86", -- $0282d
          10286 => x"86", -- $0282e
          10287 => x"85", -- $0282f
          10288 => x"83", -- $02830
          10289 => x"82", -- $02831
          10290 => x"81", -- $02832
          10291 => x"80", -- $02833
          10292 => x"80", -- $02834
          10293 => x"7f", -- $02835
          10294 => x"7f", -- $02836
          10295 => x"80", -- $02837
          10296 => x"80", -- $02838
          10297 => x"80", -- $02839
          10298 => x"80", -- $0283a
          10299 => x"80", -- $0283b
          10300 => x"81", -- $0283c
          10301 => x"83", -- $0283d
          10302 => x"83", -- $0283e
          10303 => x"82", -- $0283f
          10304 => x"81", -- $02840
          10305 => x"80", -- $02841
          10306 => x"7f", -- $02842
          10307 => x"7e", -- $02843
          10308 => x"7d", -- $02844
          10309 => x"7b", -- $02845
          10310 => x"7a", -- $02846
          10311 => x"79", -- $02847
          10312 => x"7a", -- $02848
          10313 => x"7a", -- $02849
          10314 => x"7b", -- $0284a
          10315 => x"7b", -- $0284b
          10316 => x"7c", -- $0284c
          10317 => x"7e", -- $0284d
          10318 => x"80", -- $0284e
          10319 => x"80", -- $0284f
          10320 => x"7e", -- $02850
          10321 => x"7d", -- $02851
          10322 => x"7c", -- $02852
          10323 => x"7d", -- $02853
          10324 => x"7b", -- $02854
          10325 => x"7a", -- $02855
          10326 => x"79", -- $02856
          10327 => x"78", -- $02857
          10328 => x"79", -- $02858
          10329 => x"7a", -- $02859
          10330 => x"7b", -- $0285a
          10331 => x"7b", -- $0285b
          10332 => x"7b", -- $0285c
          10333 => x"7e", -- $0285d
          10334 => x"80", -- $0285e
          10335 => x"81", -- $0285f
          10336 => x"83", -- $02860
          10337 => x"84", -- $02861
          10338 => x"85", -- $02862
          10339 => x"86", -- $02863
          10340 => x"87", -- $02864
          10341 => x"88", -- $02865
          10342 => x"88", -- $02866
          10343 => x"89", -- $02867
          10344 => x"86", -- $02868
          10345 => x"7b", -- $02869
          10346 => x"7b", -- $0286a
          10347 => x"80", -- $0286b
          10348 => x"7e", -- $0286c
          10349 => x"80", -- $0286d
          10350 => x"7e", -- $0286e
          10351 => x"7c", -- $0286f
          10352 => x"7e", -- $02870
          10353 => x"81", -- $02871
          10354 => x"85", -- $02872
          10355 => x"82", -- $02873
          10356 => x"7f", -- $02874
          10357 => x"7d", -- $02875
          10358 => x"7d", -- $02876
          10359 => x"7d", -- $02877
          10360 => x"7e", -- $02878
          10361 => x"7b", -- $02879
          10362 => x"76", -- $0287a
          10363 => x"79", -- $0287b
          10364 => x"7d", -- $0287c
          10365 => x"80", -- $0287d
          10366 => x"81", -- $0287e
          10367 => x"80", -- $0287f
          10368 => x"80", -- $02880
          10369 => x"81", -- $02881
          10370 => x"86", -- $02882
          10371 => x"88", -- $02883
          10372 => x"84", -- $02884
          10373 => x"80", -- $02885
          10374 => x"7e", -- $02886
          10375 => x"7d", -- $02887
          10376 => x"7d", -- $02888
          10377 => x"7b", -- $02889
          10378 => x"77", -- $0288a
          10379 => x"74", -- $0288b
          10380 => x"75", -- $0288c
          10381 => x"78", -- $0288d
          10382 => x"7b", -- $0288e
          10383 => x"7c", -- $0288f
          10384 => x"7c", -- $02890
          10385 => x"7d", -- $02891
          10386 => x"80", -- $02892
          10387 => x"84", -- $02893
          10388 => x"85", -- $02894
          10389 => x"83", -- $02895
          10390 => x"80", -- $02896
          10391 => x"7f", -- $02897
          10392 => x"7f", -- $02898
          10393 => x"7d", -- $02899
          10394 => x"7a", -- $0289a
          10395 => x"78", -- $0289b
          10396 => x"77", -- $0289c
          10397 => x"77", -- $0289d
          10398 => x"79", -- $0289e
          10399 => x"7c", -- $0289f
          10400 => x"7e", -- $028a0
          10401 => x"7f", -- $028a1
          10402 => x"80", -- $028a2
          10403 => x"84", -- $028a3
          10404 => x"85", -- $028a4
          10405 => x"86", -- $028a5
          10406 => x"84", -- $028a6
          10407 => x"83", -- $028a7
          10408 => x"81", -- $028a8
          10409 => x"81", -- $028a9
          10410 => x"80", -- $028aa
          10411 => x"7e", -- $028ab
          10412 => x"7d", -- $028ac
          10413 => x"7c", -- $028ad
          10414 => x"7d", -- $028ae
          10415 => x"7e", -- $028af
          10416 => x"7f", -- $028b0
          10417 => x"80", -- $028b1
          10418 => x"80", -- $028b2
          10419 => x"82", -- $028b3
          10420 => x"83", -- $028b4
          10421 => x"83", -- $028b5
          10422 => x"83", -- $028b6
          10423 => x"81", -- $028b7
          10424 => x"80", -- $028b8
          10425 => x"80", -- $028b9
          10426 => x"7f", -- $028ba
          10427 => x"7d", -- $028bb
          10428 => x"7c", -- $028bc
          10429 => x"7c", -- $028bd
          10430 => x"7c", -- $028be
          10431 => x"7d", -- $028bf
          10432 => x"7e", -- $028c0
          10433 => x"7e", -- $028c1
          10434 => x"80", -- $028c2
          10435 => x"80", -- $028c3
          10436 => x"81", -- $028c4
          10437 => x"81", -- $028c5
          10438 => x"82", -- $028c6
          10439 => x"81", -- $028c7
          10440 => x"80", -- $028c8
          10441 => x"80", -- $028c9
          10442 => x"7e", -- $028ca
          10443 => x"7e", -- $028cb
          10444 => x"7e", -- $028cc
          10445 => x"7d", -- $028cd
          10446 => x"7c", -- $028ce
          10447 => x"7c", -- $028cf
          10448 => x"7e", -- $028d0
          10449 => x"7f", -- $028d1
          10450 => x"80", -- $028d2
          10451 => x"80", -- $028d3
          10452 => x"80", -- $028d4
          10453 => x"81", -- $028d5
          10454 => x"81", -- $028d6
          10455 => x"82", -- $028d7
          10456 => x"80", -- $028d8
          10457 => x"80", -- $028d9
          10458 => x"7f", -- $028da
          10459 => x"7e", -- $028db
          10460 => x"7f", -- $028dc
          10461 => x"7e", -- $028dd
          10462 => x"7d", -- $028de
          10463 => x"7c", -- $028df
          10464 => x"7d", -- $028e0
          10465 => x"80", -- $028e1
          10466 => x"80", -- $028e2
          10467 => x"81", -- $028e3
          10468 => x"82", -- $028e4
          10469 => x"82", -- $028e5
          10470 => x"84", -- $028e6
          10471 => x"85", -- $028e7
          10472 => x"85", -- $028e8
          10473 => x"84", -- $028e9
          10474 => x"82", -- $028ea
          10475 => x"81", -- $028eb
          10476 => x"81", -- $028ec
          10477 => x"80", -- $028ed
          10478 => x"80", -- $028ee
          10479 => x"80", -- $028ef
          10480 => x"80", -- $028f0
          10481 => x"80", -- $028f1
          10482 => x"80", -- $028f2
          10483 => x"80", -- $028f3
          10484 => x"80", -- $028f4
          10485 => x"80", -- $028f5
          10486 => x"80", -- $028f6
          10487 => x"81", -- $028f7
          10488 => x"81", -- $028f8
          10489 => x"81", -- $028f9
          10490 => x"80", -- $028fa
          10491 => x"80", -- $028fb
          10492 => x"80", -- $028fc
          10493 => x"80", -- $028fd
          10494 => x"80", -- $028fe
          10495 => x"80", -- $028ff
          10496 => x"80", -- $02900
          10497 => x"80", -- $02901
          10498 => x"81", -- $02902
          10499 => x"81", -- $02903
          10500 => x"81", -- $02904
          10501 => x"80", -- $02905
          10502 => x"80", -- $02906
          10503 => x"80", -- $02907
          10504 => x"81", -- $02908
          10505 => x"80", -- $02909
          10506 => x"80", -- $0290a
          10507 => x"7f", -- $0290b
          10508 => x"7f", -- $0290c
          10509 => x"7f", -- $0290d
          10510 => x"7f", -- $0290e
          10511 => x"7e", -- $0290f
          10512 => x"7e", -- $02910
          10513 => x"7e", -- $02911
          10514 => x"7f", -- $02912
          10515 => x"7f", -- $02913
          10516 => x"80", -- $02914
          10517 => x"80", -- $02915
          10518 => x"80", -- $02916
          10519 => x"80", -- $02917
          10520 => x"81", -- $02918
          10521 => x"82", -- $02919
          10522 => x"82", -- $0291a
          10523 => x"82", -- $0291b
          10524 => x"82", -- $0291c
          10525 => x"83", -- $0291d
          10526 => x"83", -- $0291e
          10527 => x"82", -- $0291f
          10528 => x"82", -- $02920
          10529 => x"82", -- $02921
          10530 => x"82", -- $02922
          10531 => x"82", -- $02923
          10532 => x"82", -- $02924
          10533 => x"82", -- $02925
          10534 => x"82", -- $02926
          10535 => x"81", -- $02927
          10536 => x"82", -- $02928
          10537 => x"82", -- $02929
          10538 => x"81", -- $0292a
          10539 => x"80", -- $0292b
          10540 => x"80", -- $0292c
          10541 => x"80", -- $0292d
          10542 => x"7f", -- $0292e
          10543 => x"7f", -- $0292f
          10544 => x"80", -- $02930
          10545 => x"7f", -- $02931
          10546 => x"80", -- $02932
          10547 => x"80", -- $02933
          10548 => x"80", -- $02934
          10549 => x"81", -- $02935
          10550 => x"80", -- $02936
          10551 => x"81", -- $02937
          10552 => x"80", -- $02938
          10553 => x"80", -- $02939
          10554 => x"81", -- $0293a
          10555 => x"81", -- $0293b
          10556 => x"81", -- $0293c
          10557 => x"82", -- $0293d
          10558 => x"82", -- $0293e
          10559 => x"84", -- $0293f
          10560 => x"87", -- $02940
          10561 => x"8a", -- $02941
          10562 => x"80", -- $02942
          10563 => x"7b", -- $02943
          10564 => x"83", -- $02944
          10565 => x"81", -- $02945
          10566 => x"83", -- $02946
          10567 => x"81", -- $02947
          10568 => x"7d", -- $02948
          10569 => x"7f", -- $02949
          10570 => x"80", -- $0294a
          10571 => x"85", -- $0294b
          10572 => x"81", -- $0294c
          10573 => x"7d", -- $0294d
          10574 => x"7c", -- $0294e
          10575 => x"7e", -- $0294f
          10576 => x"7f", -- $02950
          10577 => x"7f", -- $02951
          10578 => x"7c", -- $02952
          10579 => x"78", -- $02953
          10580 => x"7c", -- $02954
          10581 => x"81", -- $02955
          10582 => x"84", -- $02956
          10583 => x"83", -- $02957
          10584 => x"80", -- $02958
          10585 => x"82", -- $02959
          10586 => x"84", -- $0295a
          10587 => x"87", -- $0295b
          10588 => x"87", -- $0295c
          10589 => x"81", -- $0295d
          10590 => x"7f", -- $0295e
          10591 => x"80", -- $0295f
          10592 => x"81", -- $02960
          10593 => x"80", -- $02961
          10594 => x"7e", -- $02962
          10595 => x"7b", -- $02963
          10596 => x"7c", -- $02964
          10597 => x"80", -- $02965
          10598 => x"82", -- $02966
          10599 => x"81", -- $02967
          10600 => x"80", -- $02968
          10601 => x"82", -- $02969
          10602 => x"85", -- $0296a
          10603 => x"87", -- $0296b
          10604 => x"87", -- $0296c
          10605 => x"83", -- $0296d
          10606 => x"82", -- $0296e
          10607 => x"82", -- $0296f
          10608 => x"83", -- $02970
          10609 => x"80", -- $02971
          10610 => x"7e", -- $02972
          10611 => x"7b", -- $02973
          10612 => x"7b", -- $02974
          10613 => x"7d", -- $02975
          10614 => x"7e", -- $02976
          10615 => x"7e", -- $02977
          10616 => x"7e", -- $02978
          10617 => x"7f", -- $02979
          10618 => x"82", -- $0297a
          10619 => x"84", -- $0297b
          10620 => x"84", -- $0297c
          10621 => x"83", -- $0297d
          10622 => x"81", -- $0297e
          10623 => x"82", -- $0297f
          10624 => x"83", -- $02980
          10625 => x"80", -- $02981
          10626 => x"80", -- $02982
          10627 => x"7d", -- $02983
          10628 => x"7c", -- $02984
          10629 => x"7e", -- $02985
          10630 => x"7e", -- $02986
          10631 => x"7e", -- $02987
          10632 => x"7e", -- $02988
          10633 => x"80", -- $02989
          10634 => x"81", -- $0298a
          10635 => x"83", -- $0298b
          10636 => x"83", -- $0298c
          10637 => x"83", -- $0298d
          10638 => x"83", -- $0298e
          10639 => x"84", -- $0298f
          10640 => x"84", -- $02990
          10641 => x"81", -- $02991
          10642 => x"80", -- $02992
          10643 => x"80", -- $02993
          10644 => x"7f", -- $02994
          10645 => x"7f", -- $02995
          10646 => x"80", -- $02996
          10647 => x"80", -- $02997
          10648 => x"80", -- $02998
          10649 => x"82", -- $02999
          10650 => x"82", -- $0299a
          10651 => x"83", -- $0299b
          10652 => x"85", -- $0299c
          10653 => x"85", -- $0299d
          10654 => x"85", -- $0299e
          10655 => x"85", -- $0299f
          10656 => x"84", -- $029a0
          10657 => x"82", -- $029a1
          10658 => x"81", -- $029a2
          10659 => x"80", -- $029a3
          10660 => x"7f", -- $029a4
          10661 => x"7f", -- $029a5
          10662 => x"7e", -- $029a6
          10663 => x"7d", -- $029a7
          10664 => x"7e", -- $029a8
          10665 => x"7f", -- $029a9
          10666 => x"80", -- $029aa
          10667 => x"80", -- $029ab
          10668 => x"82", -- $029ac
          10669 => x"83", -- $029ad
          10670 => x"84", -- $029ae
          10671 => x"85", -- $029af
          10672 => x"85", -- $029b0
          10673 => x"83", -- $029b1
          10674 => x"82", -- $029b2
          10675 => x"82", -- $029b3
          10676 => x"80", -- $029b4
          10677 => x"80", -- $029b5
          10678 => x"7f", -- $029b6
          10679 => x"7e", -- $029b7
          10680 => x"7e", -- $029b8
          10681 => x"7f", -- $029b9
          10682 => x"80", -- $029ba
          10683 => x"80", -- $029bb
          10684 => x"82", -- $029bc
          10685 => x"83", -- $029bd
          10686 => x"84", -- $029be
          10687 => x"85", -- $029bf
          10688 => x"84", -- $029c0
          10689 => x"84", -- $029c1
          10690 => x"83", -- $029c2
          10691 => x"82", -- $029c3
          10692 => x"80", -- $029c4
          10693 => x"80", -- $029c5
          10694 => x"7f", -- $029c6
          10695 => x"7e", -- $029c7
          10696 => x"7d", -- $029c8
          10697 => x"7d", -- $029c9
          10698 => x"7e", -- $029ca
          10699 => x"7f", -- $029cb
          10700 => x"80", -- $029cc
          10701 => x"81", -- $029cd
          10702 => x"81", -- $029ce
          10703 => x"82", -- $029cf
          10704 => x"83", -- $029d0
          10705 => x"83", -- $029d1
          10706 => x"83", -- $029d2
          10707 => x"82", -- $029d3
          10708 => x"82", -- $029d4
          10709 => x"81", -- $029d5
          10710 => x"81", -- $029d6
          10711 => x"80", -- $029d7
          10712 => x"80", -- $029d8
          10713 => x"80", -- $029d9
          10714 => x"80", -- $029da
          10715 => x"80", -- $029db
          10716 => x"81", -- $029dc
          10717 => x"82", -- $029dd
          10718 => x"81", -- $029de
          10719 => x"83", -- $029df
          10720 => x"83", -- $029e0
          10721 => x"84", -- $029e1
          10722 => x"84", -- $029e2
          10723 => x"83", -- $029e3
          10724 => x"83", -- $029e4
          10725 => x"82", -- $029e5
          10726 => x"81", -- $029e6
          10727 => x"80", -- $029e7
          10728 => x"80", -- $029e8
          10729 => x"80", -- $029e9
          10730 => x"7f", -- $029ea
          10731 => x"80", -- $029eb
          10732 => x"7f", -- $029ec
          10733 => x"7f", -- $029ed
          10734 => x"80", -- $029ee
          10735 => x"80", -- $029ef
          10736 => x"80", -- $029f0
          10737 => x"81", -- $029f1
          10738 => x"81", -- $029f2
          10739 => x"81", -- $029f3
          10740 => x"82", -- $029f4
          10741 => x"82", -- $029f5
          10742 => x"81", -- $029f6
          10743 => x"81", -- $029f7
          10744 => x"80", -- $029f8
          10745 => x"80", -- $029f9
          10746 => x"80", -- $029fa
          10747 => x"80", -- $029fb
          10748 => x"80", -- $029fc
          10749 => x"80", -- $029fd
          10750 => x"80", -- $029fe
          10751 => x"81", -- $029ff
          10752 => x"81", -- $02a00
          10753 => x"81", -- $02a01
          10754 => x"80", -- $02a02
          10755 => x"81", -- $02a03
          10756 => x"83", -- $02a04
          10757 => x"81", -- $02a05
          10758 => x"82", -- $02a06
          10759 => x"81", -- $02a07
          10760 => x"82", -- $02a08
          10761 => x"82", -- $02a09
          10762 => x"81", -- $02a0a
          10763 => x"80", -- $02a0b
          10764 => x"80", -- $02a0c
          10765 => x"80", -- $02a0d
          10766 => x"80", -- $02a0e
          10767 => x"80", -- $02a0f
          10768 => x"7f", -- $02a10
          10769 => x"80", -- $02a11
          10770 => x"80", -- $02a12
          10771 => x"80", -- $02a13
          10772 => x"80", -- $02a14
          10773 => x"80", -- $02a15
          10774 => x"80", -- $02a16
          10775 => x"80", -- $02a17
          10776 => x"81", -- $02a18
          10777 => x"80", -- $02a19
          10778 => x"80", -- $02a1a
          10779 => x"80", -- $02a1b
          10780 => x"80", -- $02a1c
          10781 => x"80", -- $02a1d
          10782 => x"7f", -- $02a1e
          10783 => x"7f", -- $02a1f
          10784 => x"7f", -- $02a20
          10785 => x"7f", -- $02a21
          10786 => x"7f", -- $02a22
          10787 => x"7f", -- $02a23
          10788 => x"80", -- $02a24
          10789 => x"80", -- $02a25
          10790 => x"81", -- $02a26
          10791 => x"81", -- $02a27
          10792 => x"82", -- $02a28
          10793 => x"82", -- $02a29
          10794 => x"83", -- $02a2a
          10795 => x"83", -- $02a2b
          10796 => x"82", -- $02a2c
          10797 => x"82", -- $02a2d
          10798 => x"81", -- $02a2e
          10799 => x"80", -- $02a2f
          10800 => x"80", -- $02a30
          10801 => x"80", -- $02a31
          10802 => x"7e", -- $02a32
          10803 => x"7e", -- $02a33
          10804 => x"7e", -- $02a34
          10805 => x"7e", -- $02a35
          10806 => x"7f", -- $02a36
          10807 => x"7f", -- $02a37
          10808 => x"80", -- $02a38
          10809 => x"80", -- $02a39
          10810 => x"81", -- $02a3a
          10811 => x"81", -- $02a3b
          10812 => x"80", -- $02a3c
          10813 => x"81", -- $02a3d
          10814 => x"81", -- $02a3e
          10815 => x"80", -- $02a3f
          10816 => x"80", -- $02a40
          10817 => x"80", -- $02a41
          10818 => x"80", -- $02a42
          10819 => x"7f", -- $02a43
          10820 => x"7f", -- $02a44
          10821 => x"7f", -- $02a45
          10822 => x"7e", -- $02a46
          10823 => x"80", -- $02a47
          10824 => x"80", -- $02a48
          10825 => x"80", -- $02a49
          10826 => x"80", -- $02a4a
          10827 => x"80", -- $02a4b
          10828 => x"82", -- $02a4c
          10829 => x"82", -- $02a4d
          10830 => x"81", -- $02a4e
          10831 => x"81", -- $02a4f
          10832 => x"81", -- $02a50
          10833 => x"81", -- $02a51
          10834 => x"81", -- $02a52
          10835 => x"80", -- $02a53
          10836 => x"80", -- $02a54
          10837 => x"80", -- $02a55
          10838 => x"80", -- $02a56
          10839 => x"80", -- $02a57
          10840 => x"80", -- $02a58
          10841 => x"80", -- $02a59
          10842 => x"80", -- $02a5a
          10843 => x"81", -- $02a5b
          10844 => x"81", -- $02a5c
          10845 => x"81", -- $02a5d
          10846 => x"82", -- $02a5e
          10847 => x"81", -- $02a5f
          10848 => x"81", -- $02a60
          10849 => x"80", -- $02a61
          10850 => x"80", -- $02a62
          10851 => x"80", -- $02a63
          10852 => x"80", -- $02a64
          10853 => x"7f", -- $02a65
          10854 => x"7f", -- $02a66
          10855 => x"7f", -- $02a67
          10856 => x"7f", -- $02a68
          10857 => x"7f", -- $02a69
          10858 => x"7f", -- $02a6a
          10859 => x"80", -- $02a6b
          10860 => x"80", -- $02a6c
          10861 => x"80", -- $02a6d
          10862 => x"80", -- $02a6e
          10863 => x"80", -- $02a6f
          10864 => x"80", -- $02a70
          10865 => x"81", -- $02a71
          10866 => x"81", -- $02a72
          10867 => x"80", -- $02a73
          10868 => x"80", -- $02a74
          10869 => x"80", -- $02a75
          10870 => x"80", -- $02a76
          10871 => x"80", -- $02a77
          10872 => x"80", -- $02a78
          10873 => x"7f", -- $02a79
          10874 => x"80", -- $02a7a
          10875 => x"80", -- $02a7b
          10876 => x"81", -- $02a7c
          10877 => x"80", -- $02a7d
          10878 => x"81", -- $02a7e
          10879 => x"81", -- $02a7f
          10880 => x"81", -- $02a80
          10881 => x"81", -- $02a81
          10882 => x"80", -- $02a82
          10883 => x"80", -- $02a83
          10884 => x"80", -- $02a84
          10885 => x"80", -- $02a85
          10886 => x"80", -- $02a86
          10887 => x"7f", -- $02a87
          10888 => x"7f", -- $02a88
          10889 => x"7f", -- $02a89
          10890 => x"7f", -- $02a8a
          10891 => x"7e", -- $02a8b
          10892 => x"7f", -- $02a8c
          10893 => x"80", -- $02a8d
          10894 => x"80", -- $02a8e
          10895 => x"80", -- $02a8f
          10896 => x"80", -- $02a90
          10897 => x"80", -- $02a91
          10898 => x"81", -- $02a92
          10899 => x"80", -- $02a93
          10900 => x"80", -- $02a94
          10901 => x"80", -- $02a95
          10902 => x"81", -- $02a96
          10903 => x"80", -- $02a97
          10904 => x"80", -- $02a98
          10905 => x"80", -- $02a99
          10906 => x"81", -- $02a9a
          10907 => x"82", -- $02a9b
          10908 => x"81", -- $02a9c
          10909 => x"7f", -- $02a9d
          10910 => x"80", -- $02a9e
          10911 => x"81", -- $02a9f
          10912 => x"81", -- $02aa0
          10913 => x"80", -- $02aa1
          10914 => x"80", -- $02aa2
          10915 => x"82", -- $02aa3
          10916 => x"82", -- $02aa4
          10917 => x"81", -- $02aa5
          10918 => x"80", -- $02aa6
          10919 => x"80", -- $02aa7
          10920 => x"81", -- $02aa8
          10921 => x"80", -- $02aa9
          10922 => x"7e", -- $02aaa
          10923 => x"7e", -- $02aab
          10924 => x"7e", -- $02aac
          10925 => x"7e", -- $02aad
          10926 => x"7d", -- $02aae
          10927 => x"7c", -- $02aaf
          10928 => x"7e", -- $02ab0
          10929 => x"7f", -- $02ab1
          10930 => x"7f", -- $02ab2
          10931 => x"7f", -- $02ab3
          10932 => x"7f", -- $02ab4
          10933 => x"80", -- $02ab5
          10934 => x"80", -- $02ab6
          10935 => x"80", -- $02ab7
          10936 => x"80", -- $02ab8
          10937 => x"80", -- $02ab9
          10938 => x"80", -- $02aba
          10939 => x"80", -- $02abb
          10940 => x"7f", -- $02abc
          10941 => x"7f", -- $02abd
          10942 => x"7f", -- $02abe
          10943 => x"7f", -- $02abf
          10944 => x"7e", -- $02ac0
          10945 => x"7e", -- $02ac1
          10946 => x"7f", -- $02ac2
          10947 => x"7f", -- $02ac3
          10948 => x"80", -- $02ac4
          10949 => x"80", -- $02ac5
          10950 => x"81", -- $02ac6
          10951 => x"81", -- $02ac7
          10952 => x"82", -- $02ac8
          10953 => x"82", -- $02ac9
          10954 => x"82", -- $02aca
          10955 => x"82", -- $02acb
          10956 => x"82", -- $02acc
          10957 => x"80", -- $02acd
          10958 => x"80", -- $02ace
          10959 => x"7f", -- $02acf
          10960 => x"7f", -- $02ad0
          10961 => x"7e", -- $02ad1
          10962 => x"7d", -- $02ad2
          10963 => x"7c", -- $02ad3
          10964 => x"7c", -- $02ad4
          10965 => x"7d", -- $02ad5
          10966 => x"7d", -- $02ad6
          10967 => x"7e", -- $02ad7
          10968 => x"7f", -- $02ad8
          10969 => x"80", -- $02ad9
          10970 => x"80", -- $02ada
          10971 => x"80", -- $02adb
          10972 => x"80", -- $02adc
          10973 => x"80", -- $02add
          10974 => x"80", -- $02ade
          10975 => x"80", -- $02adf
          10976 => x"80", -- $02ae0
          10977 => x"80", -- $02ae1
          10978 => x"7f", -- $02ae2
          10979 => x"7f", -- $02ae3
          10980 => x"80", -- $02ae4
          10981 => x"7f", -- $02ae5
          10982 => x"7e", -- $02ae6
          10983 => x"7f", -- $02ae7
          10984 => x"7f", -- $02ae8
          10985 => x"7f", -- $02ae9
          10986 => x"80", -- $02aea
          10987 => x"80", -- $02aeb
          10988 => x"80", -- $02aec
          10989 => x"80", -- $02aed
          10990 => x"80", -- $02aee
          10991 => x"80", -- $02aef
          10992 => x"80", -- $02af0
          10993 => x"80", -- $02af1
          10994 => x"80", -- $02af2
          10995 => x"80", -- $02af3
          10996 => x"7f", -- $02af4
          10997 => x"7f", -- $02af5
          10998 => x"7f", -- $02af6
          10999 => x"7f", -- $02af7
          11000 => x"7f", -- $02af8
          11001 => x"7e", -- $02af9
          11002 => x"7f", -- $02afa
          11003 => x"80", -- $02afb
          11004 => x"7f", -- $02afc
          11005 => x"7f", -- $02afd
          11006 => x"7f", -- $02afe
          11007 => x"80", -- $02aff
          11008 => x"7f", -- $02b00
          11009 => x"7f", -- $02b01
          11010 => x"7e", -- $02b02
          11011 => x"7f", -- $02b03
          11012 => x"7e", -- $02b04
          11013 => x"7e", -- $02b05
          11014 => x"7e", -- $02b06
          11015 => x"7e", -- $02b07
          11016 => x"7f", -- $02b08
          11017 => x"7f", -- $02b09
          11018 => x"80", -- $02b0a
          11019 => x"7f", -- $02b0b
          11020 => x"80", -- $02b0c
          11021 => x"80", -- $02b0d
          11022 => x"80", -- $02b0e
          11023 => x"80", -- $02b0f
          11024 => x"80", -- $02b10
          11025 => x"80", -- $02b11
          11026 => x"7f", -- $02b12
          11027 => x"80", -- $02b13
          11028 => x"7e", -- $02b14
          11029 => x"7f", -- $02b15
          11030 => x"7f", -- $02b16
          11031 => x"7f", -- $02b17
          11032 => x"7f", -- $02b18
          11033 => x"7f", -- $02b19
          11034 => x"7f", -- $02b1a
          11035 => x"7f", -- $02b1b
          11036 => x"80", -- $02b1c
          11037 => x"80", -- $02b1d
          11038 => x"80", -- $02b1e
          11039 => x"80", -- $02b1f
          11040 => x"80", -- $02b20
          11041 => x"80", -- $02b21
          11042 => x"7f", -- $02b22
          11043 => x"7f", -- $02b23
          11044 => x"7f", -- $02b24
          11045 => x"7f", -- $02b25
          11046 => x"7e", -- $02b26
          11047 => x"7e", -- $02b27
          11048 => x"7e", -- $02b28
          11049 => x"7d", -- $02b29
          11050 => x"7e", -- $02b2a
          11051 => x"7d", -- $02b2b
          11052 => x"7e", -- $02b2c
          11053 => x"7f", -- $02b2d
          11054 => x"7f", -- $02b2e
          11055 => x"7f", -- $02b2f
          11056 => x"80", -- $02b30
          11057 => x"80", -- $02b31
          11058 => x"80", -- $02b32
          11059 => x"80", -- $02b33
          11060 => x"81", -- $02b34
          11061 => x"80", -- $02b35
          11062 => x"80", -- $02b36
          11063 => x"7f", -- $02b37
          11064 => x"80", -- $02b38
          11065 => x"7f", -- $02b39
          11066 => x"7d", -- $02b3a
          11067 => x"7f", -- $02b3b
          11068 => x"7f", -- $02b3c
          11069 => x"7f", -- $02b3d
          11070 => x"7f", -- $02b3e
          11071 => x"7f", -- $02b3f
          11072 => x"7f", -- $02b40
          11073 => x"80", -- $02b41
          11074 => x"80", -- $02b42
          11075 => x"7f", -- $02b43
          11076 => x"80", -- $02b44
          11077 => x"80", -- $02b45
          11078 => x"80", -- $02b46
          11079 => x"7f", -- $02b47
          11080 => x"7f", -- $02b48
          11081 => x"7f", -- $02b49
          11082 => x"7e", -- $02b4a
          11083 => x"7e", -- $02b4b
          11084 => x"7e", -- $02b4c
          11085 => x"7f", -- $02b4d
          11086 => x"7e", -- $02b4e
          11087 => x"7e", -- $02b4f
          11088 => x"7f", -- $02b50
          11089 => x"7f", -- $02b51
          11090 => x"80", -- $02b52
          11091 => x"7e", -- $02b53
          11092 => x"80", -- $02b54
          11093 => x"7f", -- $02b55
          11094 => x"80", -- $02b56
          11095 => x"80", -- $02b57
          11096 => x"80", -- $02b58
          11097 => x"80", -- $02b59
          11098 => x"7f", -- $02b5a
          11099 => x"80", -- $02b5b
          11100 => x"80", -- $02b5c
          11101 => x"80", -- $02b5d
          11102 => x"7f", -- $02b5e
          11103 => x"7f", -- $02b5f
          11104 => x"80", -- $02b60
          11105 => x"80", -- $02b61
          11106 => x"7f", -- $02b62
          11107 => x"80", -- $02b63
          11108 => x"80", -- $02b64
          11109 => x"80", -- $02b65
          11110 => x"80", -- $02b66
          11111 => x"80", -- $02b67
          11112 => x"80", -- $02b68
          11113 => x"80", -- $02b69
          11114 => x"80", -- $02b6a
          11115 => x"80", -- $02b6b
          11116 => x"80", -- $02b6c
          11117 => x"80", -- $02b6d
          11118 => x"7e", -- $02b6e
          11119 => x"7f", -- $02b6f
          11120 => x"7f", -- $02b70
          11121 => x"7f", -- $02b71
          11122 => x"7e", -- $02b72
          11123 => x"7f", -- $02b73
          11124 => x"80", -- $02b74
          11125 => x"7e", -- $02b75
          11126 => x"7f", -- $02b76
          11127 => x"7f", -- $02b77
          11128 => x"80", -- $02b78
          11129 => x"80", -- $02b79
          11130 => x"7f", -- $02b7a
          11131 => x"80", -- $02b7b
          11132 => x"80", -- $02b7c
          11133 => x"80", -- $02b7d
          11134 => x"7f", -- $02b7e
          11135 => x"80", -- $02b7f
          11136 => x"80", -- $02b80
          11137 => x"80", -- $02b81
          11138 => x"80", -- $02b82
          11139 => x"80", -- $02b83
          11140 => x"80", -- $02b84
          11141 => x"80", -- $02b85
          11142 => x"80", -- $02b86
          11143 => x"80", -- $02b87
          11144 => x"80", -- $02b88
          11145 => x"80", -- $02b89
          11146 => x"80", -- $02b8a
          11147 => x"80", -- $02b8b
          11148 => x"80", -- $02b8c
          11149 => x"80", -- $02b8d
          11150 => x"80", -- $02b8e
          11151 => x"80", -- $02b8f
          11152 => x"80", -- $02b90
          11153 => x"80", -- $02b91
          11154 => x"7f", -- $02b92
          11155 => x"80", -- $02b93
          11156 => x"7f", -- $02b94
          11157 => x"7f", -- $02b95
          11158 => x"80", -- $02b96
          11159 => x"80", -- $02b97
          11160 => x"80", -- $02b98
          11161 => x"80", -- $02b99
          11162 => x"80", -- $02b9a
          11163 => x"80", -- $02b9b
          11164 => x"80", -- $02b9c
          11165 => x"80", -- $02b9d
          11166 => x"80", -- $02b9e
          11167 => x"80", -- $02b9f
          11168 => x"80", -- $02ba0
          11169 => x"7e", -- $02ba1
          11170 => x"80", -- $02ba2
          11171 => x"80", -- $02ba3
          11172 => x"7f", -- $02ba4
          11173 => x"80", -- $02ba5
          11174 => x"80", -- $02ba6
          11175 => x"80", -- $02ba7
          11176 => x"80", -- $02ba8
          11177 => x"80", -- $02ba9
          11178 => x"80", -- $02baa
          11179 => x"80", -- $02bab
          11180 => x"80", -- $02bac
          11181 => x"80", -- $02bad
          11182 => x"80", -- $02bae
          11183 => x"80", -- $02baf
          11184 => x"80", -- $02bb0
          11185 => x"80", -- $02bb1
          11186 => x"80", -- $02bb2
          11187 => x"80", -- $02bb3
          11188 => x"80", -- $02bb4
          11189 => x"80", -- $02bb5
          11190 => x"80", -- $02bb6
          11191 => x"80", -- $02bb7
          11192 => x"7f", -- $02bb8
          11193 => x"80", -- $02bb9
          11194 => x"7f", -- $02bba
          11195 => x"80", -- $02bbb
          11196 => x"7f", -- $02bbc
          11197 => x"7f", -- $02bbd
          11198 => x"80", -- $02bbe
          11199 => x"80", -- $02bbf
          11200 => x"80", -- $02bc0
          11201 => x"7f", -- $02bc1
          11202 => x"80", -- $02bc2
          11203 => x"80", -- $02bc3
          11204 => x"7f", -- $02bc4
          11205 => x"80", -- $02bc5
          11206 => x"7f", -- $02bc6
          11207 => x"80", -- $02bc7
          11208 => x"80", -- $02bc8
          11209 => x"80", -- $02bc9
          11210 => x"80", -- $02bca
          11211 => x"80", -- $02bcb
          11212 => x"80", -- $02bcc
          11213 => x"80", -- $02bcd
          11214 => x"80", -- $02bce
          11215 => x"80", -- $02bcf
          11216 => x"80", -- $02bd0
          11217 => x"80", -- $02bd1
          11218 => x"80", -- $02bd2
          11219 => x"80", -- $02bd3
          11220 => x"80", -- $02bd4
          11221 => x"80", -- $02bd5
          11222 => x"80", -- $02bd6
          11223 => x"80", -- $02bd7
          11224 => x"80", -- $02bd8
          11225 => x"80", -- $02bd9
          11226 => x"80", -- $02bda
          11227 => x"80", -- $02bdb
          11228 => x"80", -- $02bdc
          11229 => x"80", -- $02bdd
          11230 => x"80", -- $02bde
          11231 => x"80", -- $02bdf
          11232 => x"80", -- $02be0
          11233 => x"80", -- $02be1
          11234 => x"80", -- $02be2
          11235 => x"7f", -- $02be3
          11236 => x"7f", -- $02be4
          11237 => x"80", -- $02be5
          11238 => x"80", -- $02be6
          11239 => x"80", -- $02be7
          11240 => x"7f", -- $02be8
          11241 => x"80", -- $02be9
          11242 => x"7f", -- $02bea
          11243 => x"80", -- $02beb
          11244 => x"80", -- $02bec
          11245 => x"80", -- $02bed
          11246 => x"80", -- $02bee
          11247 => x"80", -- $02bef
          11248 => x"80", -- $02bf0
          11249 => x"80", -- $02bf1
          11250 => x"80", -- $02bf2
          11251 => x"80", -- $02bf3
          11252 => x"80", -- $02bf4
          11253 => x"80", -- $02bf5
          11254 => x"80", -- $02bf6
          11255 => x"80", -- $02bf7
          11256 => x"80", -- $02bf8
          11257 => x"80", -- $02bf9
          11258 => x"80", -- $02bfa
          11259 => x"80", -- $02bfb
          11260 => x"80", -- $02bfc
          11261 => x"80", -- $02bfd
          11262 => x"80", -- $02bfe
          11263 => x"80", -- $02bff
          11264 => x"80", -- $02c00
          11265 => x"80", -- $02c01
          11266 => x"80", -- $02c02
          11267 => x"81", -- $02c03
          11268 => x"80", -- $02c04
          11269 => x"80", -- $02c05
          11270 => x"80", -- $02c06
          11271 => x"81", -- $02c07
          11272 => x"80", -- $02c08
          11273 => x"80", -- $02c09
          11274 => x"80", -- $02c0a
          11275 => x"80", -- $02c0b
          11276 => x"80", -- $02c0c
          11277 => x"80", -- $02c0d
          11278 => x"80", -- $02c0e
          11279 => x"80", -- $02c0f
          11280 => x"80", -- $02c10
          11281 => x"80", -- $02c11
          11282 => x"80", -- $02c12
          11283 => x"80", -- $02c13
          11284 => x"80", -- $02c14
          11285 => x"80", -- $02c15
          11286 => x"80", -- $02c16
          11287 => x"80", -- $02c17
          11288 => x"80", -- $02c18
          11289 => x"81", -- $02c19
          11290 => x"81", -- $02c1a
          11291 => x"81", -- $02c1b
          11292 => x"81", -- $02c1c
          11293 => x"81", -- $02c1d
          11294 => x"81", -- $02c1e
          11295 => x"81", -- $02c1f
          11296 => x"81", -- $02c20
          11297 => x"81", -- $02c21
          11298 => x"81", -- $02c22
          11299 => x"81", -- $02c23
          11300 => x"81", -- $02c24
          11301 => x"81", -- $02c25
          11302 => x"81", -- $02c26
          11303 => x"81", -- $02c27
          11304 => x"81", -- $02c28
          11305 => x"81", -- $02c29
          11306 => x"81", -- $02c2a
          11307 => x"81", -- $02c2b
          11308 => x"81", -- $02c2c
          11309 => x"81", -- $02c2d
          11310 => x"81", -- $02c2e
          11311 => x"81", -- $02c2f
          11312 => x"81", -- $02c30
          11313 => x"81", -- $02c31
          11314 => x"81", -- $02c32
          11315 => x"81", -- $02c33
          11316 => x"81", -- $02c34
          11317 => x"81", -- $02c35
          11318 => x"81", -- $02c36
          11319 => x"81", -- $02c37
          11320 => x"81", -- $02c38
          11321 => x"81", -- $02c39
          11322 => x"81", -- $02c3a
          11323 => x"81", -- $02c3b
          11324 => x"81", -- $02c3c
          11325 => x"81", -- $02c3d
          11326 => x"82", -- $02c3e
          11327 => x"81", -- $02c3f
          11328 => x"82", -- $02c40
          11329 => x"82", -- $02c41
          11330 => x"81", -- $02c42
          11331 => x"82", -- $02c43
          11332 => x"82", -- $02c44
          11333 => x"82", -- $02c45
          11334 => x"81", -- $02c46
          11335 => x"81", -- $02c47
          11336 => x"81", -- $02c48
          11337 => x"80", -- $02c49
          11338 => x"80", -- $02c4a
          11339 => x"80", -- $02c4b
          11340 => x"80", -- $02c4c
          11341 => x"7f", -- $02c4d
          11342 => x"80", -- $02c4e
          11343 => x"80", -- $02c4f
          11344 => x"7f", -- $02c50
          11345 => x"7f", -- $02c51
          11346 => x"80", -- $02c52
          11347 => x"80", -- $02c53
          11348 => x"80", -- $02c54
          11349 => x"80", -- $02c55
          11350 => x"80", -- $02c56
          11351 => x"80", -- $02c57
          11352 => x"81", -- $02c58
          11353 => x"82", -- $02c59
          11354 => x"82", -- $02c5a
          11355 => x"83", -- $02c5b
          11356 => x"84", -- $02c5c
          11357 => x"85", -- $02c5d
          11358 => x"85", -- $02c5e
          11359 => x"86", -- $02c5f
          11360 => x"86", -- $02c60
          11361 => x"87", -- $02c61
          11362 => x"85", -- $02c62
          11363 => x"82", -- $02c63
          11364 => x"87", -- $02c64
          11365 => x"85", -- $02c65
          11366 => x"80", -- $02c66
          11367 => x"83", -- $02c67
          11368 => x"82", -- $02c68
          11369 => x"80", -- $02c69
          11370 => x"7f", -- $02c6a
          11371 => x"80", -- $02c6b
          11372 => x"81", -- $02c6c
          11373 => x"7e", -- $02c6d
          11374 => x"7d", -- $02c6e
          11375 => x"7f", -- $02c6f
          11376 => x"80", -- $02c70
          11377 => x"7d", -- $02c71
          11378 => x"7e", -- $02c72
          11379 => x"80", -- $02c73
          11380 => x"80", -- $02c74
          11381 => x"7f", -- $02c75
          11382 => x"80", -- $02c76
          11383 => x"82", -- $02c77
          11384 => x"81", -- $02c78
          11385 => x"80", -- $02c79
          11386 => x"81", -- $02c7a
          11387 => x"83", -- $02c7b
          11388 => x"82", -- $02c7c
          11389 => x"81", -- $02c7d
          11390 => x"82", -- $02c7e
          11391 => x"83", -- $02c7f
          11392 => x"81", -- $02c80
          11393 => x"80", -- $02c81
          11394 => x"81", -- $02c82
          11395 => x"80", -- $02c83
          11396 => x"80", -- $02c84
          11397 => x"80", -- $02c85
          11398 => x"80", -- $02c86
          11399 => x"7f", -- $02c87
          11400 => x"7e", -- $02c88
          11401 => x"7f", -- $02c89
          11402 => x"7f", -- $02c8a
          11403 => x"7f", -- $02c8b
          11404 => x"80", -- $02c8c
          11405 => x"80", -- $02c8d
          11406 => x"80", -- $02c8e
          11407 => x"81", -- $02c8f
          11408 => x"81", -- $02c90
          11409 => x"82", -- $02c91
          11410 => x"83", -- $02c92
          11411 => x"82", -- $02c93
          11412 => x"83", -- $02c94
          11413 => x"82", -- $02c95
          11414 => x"82", -- $02c96
          11415 => x"81", -- $02c97
          11416 => x"80", -- $02c98
          11417 => x"81", -- $02c99
          11418 => x"80", -- $02c9a
          11419 => x"80", -- $02c9b
          11420 => x"80", -- $02c9c
          11421 => x"80", -- $02c9d
          11422 => x"80", -- $02c9e
          11423 => x"80", -- $02c9f
          11424 => x"80", -- $02ca0
          11425 => x"81", -- $02ca1
          11426 => x"80", -- $02ca2
          11427 => x"81", -- $02ca3
          11428 => x"81", -- $02ca4
          11429 => x"82", -- $02ca5
          11430 => x"82", -- $02ca6
          11431 => x"81", -- $02ca7
          11432 => x"82", -- $02ca8
          11433 => x"82", -- $02ca9
          11434 => x"82", -- $02caa
          11435 => x"81", -- $02cab
          11436 => x"81", -- $02cac
          11437 => x"81", -- $02cad
          11438 => x"80", -- $02cae
          11439 => x"80", -- $02caf
          11440 => x"80", -- $02cb0
          11441 => x"80", -- $02cb1
          11442 => x"80", -- $02cb2
          11443 => x"81", -- $02cb3
          11444 => x"80", -- $02cb4
          11445 => x"80", -- $02cb5
          11446 => x"81", -- $02cb6
          11447 => x"81", -- $02cb7
          11448 => x"81", -- $02cb8
          11449 => x"81", -- $02cb9
          11450 => x"82", -- $02cba
          11451 => x"82", -- $02cbb
          11452 => x"81", -- $02cbc
          11453 => x"81", -- $02cbd
          11454 => x"81", -- $02cbe
          11455 => x"82", -- $02cbf
          11456 => x"81", -- $02cc0
          11457 => x"81", -- $02cc1
          11458 => x"81", -- $02cc2
          11459 => x"81", -- $02cc3
          11460 => x"80", -- $02cc4
          11461 => x"80", -- $02cc5
          11462 => x"80", -- $02cc6
          11463 => x"80", -- $02cc7
          11464 => x"80", -- $02cc8
          11465 => x"80", -- $02cc9
          11466 => x"80", -- $02cca
          11467 => x"80", -- $02ccb
          11468 => x"80", -- $02ccc
          11469 => x"81", -- $02ccd
          11470 => x"82", -- $02cce
          11471 => x"82", -- $02ccf
          11472 => x"83", -- $02cd0
          11473 => x"82", -- $02cd1
          11474 => x"84", -- $02cd2
          11475 => x"83", -- $02cd3
          11476 => x"82", -- $02cd4
          11477 => x"84", -- $02cd5
          11478 => x"82", -- $02cd6
          11479 => x"82", -- $02cd7
          11480 => x"81", -- $02cd8
          11481 => x"80", -- $02cd9
          11482 => x"80", -- $02cda
          11483 => x"7f", -- $02cdb
          11484 => x"7f", -- $02cdc
          11485 => x"7e", -- $02cdd
          11486 => x"7d", -- $02cde
          11487 => x"7d", -- $02cdf
          11488 => x"7d", -- $02ce0
          11489 => x"7d", -- $02ce1
          11490 => x"7c", -- $02ce2
          11491 => x"7d", -- $02ce3
          11492 => x"7e", -- $02ce4
          11493 => x"7d", -- $02ce5
          11494 => x"7f", -- $02ce6
          11495 => x"80", -- $02ce7
          11496 => x"80", -- $02ce8
          11497 => x"80", -- $02ce9
          11498 => x"81", -- $02cea
          11499 => x"82", -- $02ceb
          11500 => x"82", -- $02cec
          11501 => x"84", -- $02ced
          11502 => x"84", -- $02cee
          11503 => x"85", -- $02cef
          11504 => x"86", -- $02cf0
          11505 => x"86", -- $02cf1
          11506 => x"87", -- $02cf2
          11507 => x"89", -- $02cf3
          11508 => x"89", -- $02cf4
          11509 => x"82", -- $02cf5
          11510 => x"87", -- $02cf6
          11511 => x"8c", -- $02cf7
          11512 => x"80", -- $02cf8
          11513 => x"84", -- $02cf9
          11514 => x"85", -- $02cfa
          11515 => x"83", -- $02cfb
          11516 => x"82", -- $02cfc
          11517 => x"7c", -- $02cfd
          11518 => x"81", -- $02cfe
          11519 => x"81", -- $02cff
          11520 => x"79", -- $02d00
          11521 => x"7b", -- $02d01
          11522 => x"80", -- $02d02
          11523 => x"7c", -- $02d03
          11524 => x"78", -- $02d04
          11525 => x"7b", -- $02d05
          11526 => x"7c", -- $02d06
          11527 => x"7d", -- $02d07
          11528 => x"7b", -- $02d08
          11529 => x"7c", -- $02d09
          11530 => x"80", -- $02d0a
          11531 => x"80", -- $02d0b
          11532 => x"7e", -- $02d0c
          11533 => x"80", -- $02d0d
          11534 => x"83", -- $02d0e
          11535 => x"83", -- $02d0f
          11536 => x"81", -- $02d10
          11537 => x"84", -- $02d11
          11538 => x"85", -- $02d12
          11539 => x"84", -- $02d13
          11540 => x"81", -- $02d14
          11541 => x"82", -- $02d15
          11542 => x"83", -- $02d16
          11543 => x"80", -- $02d17
          11544 => x"7e", -- $02d18
          11545 => x"7f", -- $02d19
          11546 => x"7e", -- $02d1a
          11547 => x"7c", -- $02d1b
          11548 => x"7b", -- $02d1c
          11549 => x"7b", -- $02d1d
          11550 => x"7e", -- $02d1e
          11551 => x"7c", -- $02d1f
          11552 => x"7c", -- $02d20
          11553 => x"80", -- $02d21
          11554 => x"80", -- $02d22
          11555 => x"80", -- $02d23
          11556 => x"80", -- $02d24
          11557 => x"82", -- $02d25
          11558 => x"83", -- $02d26
          11559 => x"83", -- $02d27
          11560 => x"83", -- $02d28
          11561 => x"83", -- $02d29
          11562 => x"85", -- $02d2a
          11563 => x"83", -- $02d2b
          11564 => x"82", -- $02d2c
          11565 => x"83", -- $02d2d
          11566 => x"82", -- $02d2e
          11567 => x"81", -- $02d2f
          11568 => x"80", -- $02d30
          11569 => x"81", -- $02d31
          11570 => x"81", -- $02d32
          11571 => x"80", -- $02d33
          11572 => x"80", -- $02d34
          11573 => x"80", -- $02d35
          11574 => x"81", -- $02d36
          11575 => x"80", -- $02d37
          11576 => x"80", -- $02d38
          11577 => x"81", -- $02d39
          11578 => x"81", -- $02d3a
          11579 => x"80", -- $02d3b
          11580 => x"80", -- $02d3c
          11581 => x"81", -- $02d3d
          11582 => x"81", -- $02d3e
          11583 => x"80", -- $02d3f
          11584 => x"80", -- $02d40
          11585 => x"80", -- $02d41
          11586 => x"80", -- $02d42
          11587 => x"80", -- $02d43
          11588 => x"7f", -- $02d44
          11589 => x"80", -- $02d45
          11590 => x"80", -- $02d46
          11591 => x"7f", -- $02d47
          11592 => x"80", -- $02d48
          11593 => x"80", -- $02d49
          11594 => x"80", -- $02d4a
          11595 => x"80", -- $02d4b
          11596 => x"80", -- $02d4c
          11597 => x"80", -- $02d4d
          11598 => x"81", -- $02d4e
          11599 => x"80", -- $02d4f
          11600 => x"80", -- $02d50
          11601 => x"80", -- $02d51
          11602 => x"80", -- $02d52
          11603 => x"80", -- $02d53
          11604 => x"80", -- $02d54
          11605 => x"80", -- $02d55
          11606 => x"7f", -- $02d56
          11607 => x"7f", -- $02d57
          11608 => x"7e", -- $02d58
          11609 => x"7e", -- $02d59
          11610 => x"7e", -- $02d5a
          11611 => x"7e", -- $02d5b
          11612 => x"7e", -- $02d5c
          11613 => x"7f", -- $02d5d
          11614 => x"80", -- $02d5e
          11615 => x"80", -- $02d5f
          11616 => x"80", -- $02d60
          11617 => x"81", -- $02d61
          11618 => x"82", -- $02d62
          11619 => x"83", -- $02d63
          11620 => x"84", -- $02d64
          11621 => x"85", -- $02d65
          11622 => x"88", -- $02d66
          11623 => x"88", -- $02d67
          11624 => x"85", -- $02d68
          11625 => x"85", -- $02d69
          11626 => x"88", -- $02d6a
          11627 => x"84", -- $02d6b
          11628 => x"84", -- $02d6c
          11629 => x"82", -- $02d6d
          11630 => x"82", -- $02d6e
          11631 => x"83", -- $02d6f
          11632 => x"7e", -- $02d70
          11633 => x"7f", -- $02d71
          11634 => x"80", -- $02d72
          11635 => x"7d", -- $02d73
          11636 => x"7c", -- $02d74
          11637 => x"7c", -- $02d75
          11638 => x"7c", -- $02d76
          11639 => x"7c", -- $02d77
          11640 => x"7b", -- $02d78
          11641 => x"7b", -- $02d79
          11642 => x"7d", -- $02d7a
          11643 => x"7e", -- $02d7b
          11644 => x"7d", -- $02d7c
          11645 => x"7d", -- $02d7d
          11646 => x"7f", -- $02d7e
          11647 => x"7f", -- $02d7f
          11648 => x"7f", -- $02d80
          11649 => x"7f", -- $02d81
          11650 => x"7f", -- $02d82
          11651 => x"80", -- $02d83
          11652 => x"80", -- $02d84
          11653 => x"7f", -- $02d85
          11654 => x"80", -- $02d86
          11655 => x"80", -- $02d87
          11656 => x"80", -- $02d88
          11657 => x"7f", -- $02d89
          11658 => x"7f", -- $02d8a
          11659 => x"80", -- $02d8b
          11660 => x"7e", -- $02d8c
          11661 => x"7c", -- $02d8d
          11662 => x"7e", -- $02d8e
          11663 => x"7e", -- $02d8f
          11664 => x"7e", -- $02d90
          11665 => x"7d", -- $02d91
          11666 => x"7d", -- $02d92
          11667 => x"80", -- $02d93
          11668 => x"80", -- $02d94
          11669 => x"80", -- $02d95
          11670 => x"81", -- $02d96
          11671 => x"83", -- $02d97
          11672 => x"82", -- $02d98
          11673 => x"83", -- $02d99
          11674 => x"83", -- $02d9a
          11675 => x"84", -- $02d9b
          11676 => x"85", -- $02d9c
          11677 => x"83", -- $02d9d
          11678 => x"83", -- $02d9e
          11679 => x"80", -- $02d9f
          11680 => x"7f", -- $02da0
          11681 => x"83", -- $02da1
          11682 => x"7f", -- $02da2
          11683 => x"7e", -- $02da3
          11684 => x"7f", -- $02da4
          11685 => x"7e", -- $02da5
          11686 => x"80", -- $02da6
          11687 => x"7c", -- $02da7
          11688 => x"7d", -- $02da8
          11689 => x"80", -- $02da9
          11690 => x"7e", -- $02daa
          11691 => x"7d", -- $02dab
          11692 => x"7d", -- $02dac
          11693 => x"7d", -- $02dad
          11694 => x"7e", -- $02dae
          11695 => x"7d", -- $02daf
          11696 => x"7b", -- $02db0
          11697 => x"7c", -- $02db1
          11698 => x"7e", -- $02db2
          11699 => x"7c", -- $02db3
          11700 => x"7c", -- $02db4
          11701 => x"7d", -- $02db5
          11702 => x"7e", -- $02db6
          11703 => x"7f", -- $02db7
          11704 => x"7e", -- $02db8
          11705 => x"80", -- $02db9
          11706 => x"80", -- $02dba
          11707 => x"80", -- $02dbb
          11708 => x"81", -- $02dbc
          11709 => x"81", -- $02dbd
          11710 => x"82", -- $02dbe
          11711 => x"82", -- $02dbf
          11712 => x"80", -- $02dc0
          11713 => x"80", -- $02dc1
          11714 => x"80", -- $02dc2
          11715 => x"7f", -- $02dc3
          11716 => x"7c", -- $02dc4
          11717 => x"7b", -- $02dc5
          11718 => x"7b", -- $02dc6
          11719 => x"7b", -- $02dc7
          11720 => x"7a", -- $02dc8
          11721 => x"7a", -- $02dc9
          11722 => x"7a", -- $02dca
          11723 => x"7c", -- $02dcb
          11724 => x"7c", -- $02dcc
          11725 => x"7c", -- $02dcd
          11726 => x"7d", -- $02dce
          11727 => x"7e", -- $02dcf
          11728 => x"7f", -- $02dd0
          11729 => x"7f", -- $02dd1
          11730 => x"80", -- $02dd2
          11731 => x"80", -- $02dd3
          11732 => x"81", -- $02dd4
          11733 => x"81", -- $02dd5
          11734 => x"82", -- $02dd6
          11735 => x"83", -- $02dd7
          11736 => x"84", -- $02dd8
          11737 => x"85", -- $02dd9
          11738 => x"82", -- $02dda
          11739 => x"84", -- $02ddb
          11740 => x"86", -- $02ddc
          11741 => x"84", -- $02ddd
          11742 => x"84", -- $02dde
          11743 => x"83", -- $02ddf
          11744 => x"83", -- $02de0
          11745 => x"84", -- $02de1
          11746 => x"81", -- $02de2
          11747 => x"80", -- $02de3
          11748 => x"81", -- $02de4
          11749 => x"80", -- $02de5
          11750 => x"7f", -- $02de6
          11751 => x"7e", -- $02de7
          11752 => x"7d", -- $02de8
          11753 => x"7d", -- $02de9
          11754 => x"7c", -- $02dea
          11755 => x"7a", -- $02deb
          11756 => x"7a", -- $02dec
          11757 => x"7c", -- $02ded
          11758 => x"7c", -- $02dee
          11759 => x"7c", -- $02def
          11760 => x"7b", -- $02df0
          11761 => x"7d", -- $02df1
          11762 => x"7e", -- $02df2
          11763 => x"7e", -- $02df3
          11764 => x"7e", -- $02df4
          11765 => x"7f", -- $02df5
          11766 => x"80", -- $02df6
          11767 => x"80", -- $02df7
          11768 => x"80", -- $02df8
          11769 => x"80", -- $02df9
          11770 => x"80", -- $02dfa
          11771 => x"80", -- $02dfb
          11772 => x"80", -- $02dfc
          11773 => x"7f", -- $02dfd
          11774 => x"80", -- $02dfe
          11775 => x"7f", -- $02dff
          11776 => x"7e", -- $02e00
          11777 => x"7d", -- $02e01
          11778 => x"7d", -- $02e02
          11779 => x"7d", -- $02e03
          11780 => x"7d", -- $02e04
          11781 => x"7c", -- $02e05
          11782 => x"7d", -- $02e06
          11783 => x"7e", -- $02e07
          11784 => x"7e", -- $02e08
          11785 => x"7f", -- $02e09
          11786 => x"7f", -- $02e0a
          11787 => x"80", -- $02e0b
          11788 => x"81", -- $02e0c
          11789 => x"81", -- $02e0d
          11790 => x"82", -- $02e0e
          11791 => x"83", -- $02e0f
          11792 => x"83", -- $02e10
          11793 => x"84", -- $02e11
          11794 => x"83", -- $02e12
          11795 => x"84", -- $02e13
          11796 => x"84", -- $02e14
          11797 => x"83", -- $02e15
          11798 => x"81", -- $02e16
          11799 => x"82", -- $02e17
          11800 => x"81", -- $02e18
          11801 => x"81", -- $02e19
          11802 => x"81", -- $02e1a
          11803 => x"80", -- $02e1b
          11804 => x"80", -- $02e1c
          11805 => x"80", -- $02e1d
          11806 => x"80", -- $02e1e
          11807 => x"80", -- $02e1f
          11808 => x"80", -- $02e20
          11809 => x"7f", -- $02e21
          11810 => x"80", -- $02e22
          11811 => x"7f", -- $02e23
          11812 => x"7f", -- $02e24
          11813 => x"7f", -- $02e25
          11814 => x"7f", -- $02e26
          11815 => x"7e", -- $02e27
          11816 => x"7e", -- $02e28
          11817 => x"7d", -- $02e29
          11818 => x"7e", -- $02e2a
          11819 => x"7d", -- $02e2b
          11820 => x"7c", -- $02e2c
          11821 => x"7e", -- $02e2d
          11822 => x"7e", -- $02e2e
          11823 => x"7f", -- $02e2f
          11824 => x"7f", -- $02e30
          11825 => x"7f", -- $02e31
          11826 => x"80", -- $02e32
          11827 => x"80", -- $02e33
          11828 => x"80", -- $02e34
          11829 => x"80", -- $02e35
          11830 => x"80", -- $02e36
          11831 => x"80", -- $02e37
          11832 => x"80", -- $02e38
          11833 => x"7e", -- $02e39
          11834 => x"7d", -- $02e3a
          11835 => x"7c", -- $02e3b
          11836 => x"7c", -- $02e3c
          11837 => x"7a", -- $02e3d
          11838 => x"7a", -- $02e3e
          11839 => x"7a", -- $02e3f
          11840 => x"7a", -- $02e40
          11841 => x"7a", -- $02e41
          11842 => x"7a", -- $02e42
          11843 => x"7b", -- $02e43
          11844 => x"7c", -- $02e44
          11845 => x"7d", -- $02e45
          11846 => x"7d", -- $02e46
          11847 => x"7f", -- $02e47
          11848 => x"80", -- $02e48
          11849 => x"80", -- $02e49
          11850 => x"81", -- $02e4a
          11851 => x"81", -- $02e4b
          11852 => x"82", -- $02e4c
          11853 => x"83", -- $02e4d
          11854 => x"83", -- $02e4e
          11855 => x"83", -- $02e4f
          11856 => x"82", -- $02e50
          11857 => x"83", -- $02e51
          11858 => x"83", -- $02e52
          11859 => x"82", -- $02e53
          11860 => x"82", -- $02e54
          11861 => x"81", -- $02e55
          11862 => x"82", -- $02e56
          11863 => x"82", -- $02e57
          11864 => x"81", -- $02e58
          11865 => x"82", -- $02e59
          11866 => x"81", -- $02e5a
          11867 => x"81", -- $02e5b
          11868 => x"81", -- $02e5c
          11869 => x"80", -- $02e5d
          11870 => x"80", -- $02e5e
          11871 => x"80", -- $02e5f
          11872 => x"80", -- $02e60
          11873 => x"80", -- $02e61
          11874 => x"80", -- $02e62
          11875 => x"7f", -- $02e63
          11876 => x"7f", -- $02e64
          11877 => x"7e", -- $02e65
          11878 => x"7d", -- $02e66
          11879 => x"7d", -- $02e67
          11880 => x"7e", -- $02e68
          11881 => x"7d", -- $02e69
          11882 => x"7c", -- $02e6a
          11883 => x"7c", -- $02e6b
          11884 => x"7c", -- $02e6c
          11885 => x"7c", -- $02e6d
          11886 => x"7b", -- $02e6e
          11887 => x"7b", -- $02e6f
          11888 => x"7b", -- $02e70
          11889 => x"7b", -- $02e71
          11890 => x"7b", -- $02e72
          11891 => x"7c", -- $02e73
          11892 => x"7b", -- $02e74
          11893 => x"7d", -- $02e75
          11894 => x"7d", -- $02e76
          11895 => x"7d", -- $02e77
          11896 => x"7d", -- $02e78
          11897 => x"7e", -- $02e79
          11898 => x"7e", -- $02e7a
          11899 => x"7e", -- $02e7b
          11900 => x"7e", -- $02e7c
          11901 => x"7f", -- $02e7d
          11902 => x"7f", -- $02e7e
          11903 => x"7f", -- $02e7f
          11904 => x"7f", -- $02e80
          11905 => x"7f", -- $02e81
          11906 => x"80", -- $02e82
          11907 => x"80", -- $02e83
          11908 => x"80", -- $02e84
          11909 => x"80", -- $02e85
          11910 => x"80", -- $02e86
          11911 => x"80", -- $02e87
          11912 => x"81", -- $02e88
          11913 => x"81", -- $02e89
          11914 => x"81", -- $02e8a
          11915 => x"82", -- $02e8b
          11916 => x"82", -- $02e8c
          11917 => x"82", -- $02e8d
          11918 => x"83", -- $02e8e
          11919 => x"83", -- $02e8f
          11920 => x"82", -- $02e90
          11921 => x"83", -- $02e91
          11922 => x"82", -- $02e92
          11923 => x"82", -- $02e93
          11924 => x"82", -- $02e94
          11925 => x"81", -- $02e95
          11926 => x"82", -- $02e96
          11927 => x"81", -- $02e97
          11928 => x"80", -- $02e98
          11929 => x"80", -- $02e99
          11930 => x"80", -- $02e9a
          11931 => x"80", -- $02e9b
          11932 => x"80", -- $02e9c
          11933 => x"80", -- $02e9d
          11934 => x"80", -- $02e9e
          11935 => x"80", -- $02e9f
          11936 => x"80", -- $02ea0
          11937 => x"80", -- $02ea1
          11938 => x"80", -- $02ea2
          11939 => x"7f", -- $02ea3
          11940 => x"7f", -- $02ea4
          11941 => x"80", -- $02ea5
          11942 => x"80", -- $02ea6
          11943 => x"7f", -- $02ea7
          11944 => x"7f", -- $02ea8
          11945 => x"7f", -- $02ea9
          11946 => x"80", -- $02eaa
          11947 => x"7f", -- $02eab
          11948 => x"7f", -- $02eac
          11949 => x"7f", -- $02ead
          11950 => x"7e", -- $02eae
          11951 => x"7e", -- $02eaf
          11952 => x"7d", -- $02eb0
          11953 => x"7d", -- $02eb1
          11954 => x"7d", -- $02eb2
          11955 => x"7c", -- $02eb3
          11956 => x"7c", -- $02eb4
          11957 => x"7c", -- $02eb5
          11958 => x"7c", -- $02eb6
          11959 => x"7c", -- $02eb7
          11960 => x"7c", -- $02eb8
          11961 => x"7c", -- $02eb9
          11962 => x"7c", -- $02eba
          11963 => x"7d", -- $02ebb
          11964 => x"7e", -- $02ebc
          11965 => x"7f", -- $02ebd
          11966 => x"7f", -- $02ebe
          11967 => x"80", -- $02ebf
          11968 => x"80", -- $02ec0
          11969 => x"81", -- $02ec1
          11970 => x"82", -- $02ec2
          11971 => x"82", -- $02ec3
          11972 => x"83", -- $02ec4
          11973 => x"83", -- $02ec5
          11974 => x"83", -- $02ec6
          11975 => x"83", -- $02ec7
          11976 => x"83", -- $02ec8
          11977 => x"83", -- $02ec9
          11978 => x"84", -- $02eca
          11979 => x"84", -- $02ecb
          11980 => x"84", -- $02ecc
          11981 => x"84", -- $02ecd
          11982 => x"84", -- $02ece
          11983 => x"84", -- $02ecf
          11984 => x"84", -- $02ed0
          11985 => x"84", -- $02ed1
          11986 => x"84", -- $02ed2
          11987 => x"84", -- $02ed3
          11988 => x"83", -- $02ed4
          11989 => x"83", -- $02ed5
          11990 => x"83", -- $02ed6
          11991 => x"82", -- $02ed7
          11992 => x"82", -- $02ed8
          11993 => x"82", -- $02ed9
          11994 => x"81", -- $02eda
          11995 => x"81", -- $02edb
          11996 => x"81", -- $02edc
          11997 => x"81", -- $02edd
          11998 => x"80", -- $02ede
          11999 => x"80", -- $02edf
          12000 => x"80", -- $02ee0
          12001 => x"80", -- $02ee1
          12002 => x"80", -- $02ee2
          12003 => x"80", -- $02ee3
          12004 => x"7f", -- $02ee4
          12005 => x"7f", -- $02ee5
          12006 => x"7f", -- $02ee6
          12007 => x"7e", -- $02ee7
          12008 => x"7e", -- $02ee8
          12009 => x"7d", -- $02ee9
          12010 => x"7d", -- $02eea
          12011 => x"7c", -- $02eeb
          12012 => x"7c", -- $02eec
          12013 => x"7c", -- $02eed
          12014 => x"7b", -- $02eee
          12015 => x"7b", -- $02eef
          12016 => x"7b", -- $02ef0
          12017 => x"7b", -- $02ef1
          12018 => x"7b", -- $02ef2
          12019 => x"7c", -- $02ef3
          12020 => x"7c", -- $02ef4
          12021 => x"7d", -- $02ef5
          12022 => x"7e", -- $02ef6
          12023 => x"7e", -- $02ef7
          12024 => x"7f", -- $02ef8
          12025 => x"7f", -- $02ef9
          12026 => x"80", -- $02efa
          12027 => x"80", -- $02efb
          12028 => x"80", -- $02efc
          12029 => x"81", -- $02efd
          12030 => x"81", -- $02efe
          12031 => x"81", -- $02eff
          12032 => x"82", -- $02f00
          12033 => x"82", -- $02f01
          12034 => x"82", -- $02f02
          12035 => x"83", -- $02f03
          12036 => x"82", -- $02f04
          12037 => x"82", -- $02f05
          12038 => x"82", -- $02f06
          12039 => x"82", -- $02f07
          12040 => x"82", -- $02f08
          12041 => x"82", -- $02f09
          12042 => x"82", -- $02f0a
          12043 => x"81", -- $02f0b
          12044 => x"82", -- $02f0c
          12045 => x"81", -- $02f0d
          12046 => x"82", -- $02f0e
          12047 => x"82", -- $02f0f
          12048 => x"82", -- $02f10
          12049 => x"83", -- $02f11
          12050 => x"82", -- $02f12
          12051 => x"83", -- $02f13
          12052 => x"83", -- $02f14
          12053 => x"83", -- $02f15
          12054 => x"83", -- $02f16
          12055 => x"83", -- $02f17
          12056 => x"82", -- $02f18
          12057 => x"82", -- $02f19
          12058 => x"83", -- $02f1a
          12059 => x"82", -- $02f1b
          12060 => x"82", -- $02f1c
          12061 => x"81", -- $02f1d
          12062 => x"81", -- $02f1e
          12063 => x"81", -- $02f1f
          12064 => x"80", -- $02f20
          12065 => x"80", -- $02f21
          12066 => x"80", -- $02f22
          12067 => x"80", -- $02f23
          12068 => x"7f", -- $02f24
          12069 => x"7f", -- $02f25
          12070 => x"7e", -- $02f26
          12071 => x"7e", -- $02f27
          12072 => x"7e", -- $02f28
          12073 => x"7d", -- $02f29
          12074 => x"7d", -- $02f2a
          12075 => x"7d", -- $02f2b
          12076 => x"7d", -- $02f2c
          12077 => x"7d", -- $02f2d
          12078 => x"7c", -- $02f2e
          12079 => x"7c", -- $02f2f
          12080 => x"7c", -- $02f30
          12081 => x"7d", -- $02f31
          12082 => x"7c", -- $02f32
          12083 => x"7d", -- $02f33
          12084 => x"7d", -- $02f34
          12085 => x"7d", -- $02f35
          12086 => x"7e", -- $02f36
          12087 => x"7e", -- $02f37
          12088 => x"7e", -- $02f38
          12089 => x"7f", -- $02f39
          12090 => x"7f", -- $02f3a
          12091 => x"80", -- $02f3b
          12092 => x"80", -- $02f3c
          12093 => x"80", -- $02f3d
          12094 => x"80", -- $02f3e
          12095 => x"80", -- $02f3f
          12096 => x"81", -- $02f40
          12097 => x"81", -- $02f41
          12098 => x"82", -- $02f42
          12099 => x"82", -- $02f43
          12100 => x"82", -- $02f44
          12101 => x"82", -- $02f45
          12102 => x"82", -- $02f46
          12103 => x"83", -- $02f47
          12104 => x"83", -- $02f48
          12105 => x"84", -- $02f49
          12106 => x"84", -- $02f4a
          12107 => x"84", -- $02f4b
          12108 => x"84", -- $02f4c
          12109 => x"85", -- $02f4d
          12110 => x"84", -- $02f4e
          12111 => x"85", -- $02f4f
          12112 => x"84", -- $02f50
          12113 => x"84", -- $02f51
          12114 => x"84", -- $02f52
          12115 => x"84", -- $02f53
          12116 => x"83", -- $02f54
          12117 => x"83", -- $02f55
          12118 => x"83", -- $02f56
          12119 => x"82", -- $02f57
          12120 => x"82", -- $02f58
          12121 => x"81", -- $02f59
          12122 => x"81", -- $02f5a
          12123 => x"81", -- $02f5b
          12124 => x"81", -- $02f5c
          12125 => x"80", -- $02f5d
          12126 => x"80", -- $02f5e
          12127 => x"80", -- $02f5f
          12128 => x"80", -- $02f60
          12129 => x"80", -- $02f61
          12130 => x"80", -- $02f62
          12131 => x"7f", -- $02f63
          12132 => x"7f", -- $02f64
          12133 => x"7f", -- $02f65
          12134 => x"7f", -- $02f66
          12135 => x"7f", -- $02f67
          12136 => x"7e", -- $02f68
          12137 => x"7f", -- $02f69
          12138 => x"7f", -- $02f6a
          12139 => x"7f", -- $02f6b
          12140 => x"7f", -- $02f6c
          12141 => x"7f", -- $02f6d
          12142 => x"80", -- $02f6e
          12143 => x"7f", -- $02f6f
          12144 => x"7f", -- $02f70
          12145 => x"80", -- $02f71
          12146 => x"80", -- $02f72
          12147 => x"80", -- $02f73
          12148 => x"80", -- $02f74
          12149 => x"80", -- $02f75
          12150 => x"80", -- $02f76
          12151 => x"80", -- $02f77
          12152 => x"80", -- $02f78
          12153 => x"80", -- $02f79
          12154 => x"80", -- $02f7a
          12155 => x"80", -- $02f7b
          12156 => x"80", -- $02f7c
          12157 => x"80", -- $02f7d
          12158 => x"81", -- $02f7e
          12159 => x"81", -- $02f7f
          12160 => x"81", -- $02f80
          12161 => x"81", -- $02f81
          12162 => x"82", -- $02f82
          12163 => x"82", -- $02f83
          12164 => x"82", -- $02f84
          12165 => x"82", -- $02f85
          12166 => x"82", -- $02f86
          12167 => x"83", -- $02f87
          12168 => x"83", -- $02f88
          12169 => x"83", -- $02f89
          12170 => x"83", -- $02f8a
          12171 => x"84", -- $02f8b
          12172 => x"84", -- $02f8c
          12173 => x"84", -- $02f8d
          12174 => x"84", -- $02f8e
          12175 => x"84", -- $02f8f
          12176 => x"85", -- $02f90
          12177 => x"84", -- $02f91
          12178 => x"84", -- $02f92
          12179 => x"84", -- $02f93
          12180 => x"84", -- $02f94
          12181 => x"84", -- $02f95
          12182 => x"83", -- $02f96
          12183 => x"83", -- $02f97
          12184 => x"83", -- $02f98
          12185 => x"83", -- $02f99
          12186 => x"82", -- $02f9a
          12187 => x"82", -- $02f9b
          12188 => x"81", -- $02f9c
          12189 => x"81", -- $02f9d
          12190 => x"81", -- $02f9e
          12191 => x"80", -- $02f9f
          12192 => x"80", -- $02fa0
          12193 => x"80", -- $02fa1
          12194 => x"80", -- $02fa2
          12195 => x"80", -- $02fa3
          12196 => x"80", -- $02fa4
          12197 => x"7f", -- $02fa5
          12198 => x"80", -- $02fa6
          12199 => x"7f", -- $02fa7
          12200 => x"7f", -- $02fa8
          12201 => x"7f", -- $02fa9
          12202 => x"7f", -- $02faa
          12203 => x"7f", -- $02fab
          12204 => x"7f", -- $02fac
          12205 => x"80", -- $02fad
          12206 => x"80", -- $02fae
          12207 => x"80", -- $02faf
          12208 => x"80", -- $02fb0
          12209 => x"80", -- $02fb1
          12210 => x"80", -- $02fb2
          12211 => x"80", -- $02fb3
          12212 => x"80", -- $02fb4
          12213 => x"81", -- $02fb5
          12214 => x"81", -- $02fb6
          12215 => x"81", -- $02fb7
          12216 => x"81", -- $02fb8
          12217 => x"81", -- $02fb9
          12218 => x"82", -- $02fba
          12219 => x"82", -- $02fbb
          12220 => x"82", -- $02fbc
          12221 => x"82", -- $02fbd
          12222 => x"82", -- $02fbe
          12223 => x"82", -- $02fbf
          12224 => x"82", -- $02fc0
          12225 => x"82", -- $02fc1
          12226 => x"82", -- $02fc2
          12227 => x"82", -- $02fc3
          12228 => x"83", -- $02fc4
          12229 => x"83", -- $02fc5
          12230 => x"83", -- $02fc6
          12231 => x"84", -- $02fc7
          12232 => x"83", -- $02fc8
          12233 => x"84", -- $02fc9
          12234 => x"84", -- $02fca
          12235 => x"84", -- $02fcb
          12236 => x"84", -- $02fcc
          12237 => x"83", -- $02fcd
          12238 => x"83", -- $02fce
          12239 => x"83", -- $02fcf
          12240 => x"83", -- $02fd0
          12241 => x"83", -- $02fd1
          12242 => x"83", -- $02fd2
          12243 => x"82", -- $02fd3
          12244 => x"82", -- $02fd4
          12245 => x"82", -- $02fd5
          12246 => x"81", -- $02fd6
          12247 => x"82", -- $02fd7
          12248 => x"81", -- $02fd8
          12249 => x"81", -- $02fd9
          12250 => x"81", -- $02fda
          12251 => x"80", -- $02fdb
          12252 => x"80", -- $02fdc
          12253 => x"80", -- $02fdd
          12254 => x"80", -- $02fde
          12255 => x"80", -- $02fdf
          12256 => x"80", -- $02fe0
          12257 => x"80", -- $02fe1
          12258 => x"80", -- $02fe2
          12259 => x"80", -- $02fe3
          12260 => x"80", -- $02fe4
          12261 => x"80", -- $02fe5
          12262 => x"80", -- $02fe6
          12263 => x"80", -- $02fe7
          12264 => x"80", -- $02fe8
          12265 => x"80", -- $02fe9
          12266 => x"80", -- $02fea
          12267 => x"80", -- $02feb
          12268 => x"80", -- $02fec
          12269 => x"80", -- $02fed
          12270 => x"80", -- $02fee
          12271 => x"80", -- $02fef
          12272 => x"80", -- $02ff0
          12273 => x"80", -- $02ff1
          12274 => x"80", -- $02ff2
          12275 => x"80", -- $02ff3
          12276 => x"80", -- $02ff4
          12277 => x"80", -- $02ff5
          12278 => x"80", -- $02ff6
          12279 => x"80", -- $02ff7
          12280 => x"80", -- $02ff8
          12281 => x"80", -- $02ff9
          12282 => x"80", -- $02ffa
          12283 => x"80", -- $02ffb
          12284 => x"81", -- $02ffc
          12285 => x"81", -- $02ffd
          12286 => x"82", -- $02ffe
          12287 => x"81", -- $02fff
          12288 => x"82", -- $03000
          12289 => x"82", -- $03001
          12290 => x"82", -- $03002
          12291 => x"82", -- $03003
          12292 => x"82", -- $03004
          12293 => x"82", -- $03005
          12294 => x"82", -- $03006
          12295 => x"83", -- $03007
          12296 => x"82", -- $03008
          12297 => x"83", -- $03009
          12298 => x"83", -- $0300a
          12299 => x"82", -- $0300b
          12300 => x"82", -- $0300c
          12301 => x"82", -- $0300d
          12302 => x"81", -- $0300e
          12303 => x"81", -- $0300f
          12304 => x"81", -- $03010
          12305 => x"81", -- $03011
          12306 => x"81", -- $03012
          12307 => x"80", -- $03013
          12308 => x"80", -- $03014
          12309 => x"80", -- $03015
          12310 => x"80", -- $03016
          12311 => x"80", -- $03017
          12312 => x"80", -- $03018
          12313 => x"80", -- $03019
          12314 => x"80", -- $0301a
          12315 => x"80", -- $0301b
          12316 => x"80", -- $0301c
          12317 => x"80", -- $0301d
          12318 => x"80", -- $0301e
          12319 => x"80", -- $0301f
          12320 => x"80", -- $03020
          12321 => x"80", -- $03021
          12322 => x"7f", -- $03022
          12323 => x"7f", -- $03023
          12324 => x"7f", -- $03024
          12325 => x"7f", -- $03025
          12326 => x"7f", -- $03026
          12327 => x"7f", -- $03027
          12328 => x"7f", -- $03028
          12329 => x"7f", -- $03029
          12330 => x"7f", -- $0302a
          12331 => x"7f", -- $0302b
          12332 => x"7f", -- $0302c
          12333 => x"80", -- $0302d
          12334 => x"80", -- $0302e
          12335 => x"80", -- $0302f
          12336 => x"80", -- $03030
          12337 => x"80", -- $03031
          12338 => x"80", -- $03032
          12339 => x"80", -- $03033
          12340 => x"80", -- $03034
          12341 => x"80", -- $03035
          12342 => x"80", -- $03036
          12343 => x"80", -- $03037
          12344 => x"81", -- $03038
          12345 => x"81", -- $03039
          12346 => x"81", -- $0303a
          12347 => x"81", -- $0303b
          12348 => x"81", -- $0303c
          12349 => x"81", -- $0303d
          12350 => x"82", -- $0303e
          12351 => x"81", -- $0303f
          12352 => x"81", -- $03040
          12353 => x"82", -- $03041
          12354 => x"81", -- $03042
          12355 => x"81", -- $03043
          12356 => x"81", -- $03044
          12357 => x"81", -- $03045
          12358 => x"81", -- $03046
          12359 => x"81", -- $03047
          12360 => x"80", -- $03048
          12361 => x"80", -- $03049
          12362 => x"81", -- $0304a
          12363 => x"80", -- $0304b
          12364 => x"81", -- $0304c
          12365 => x"80", -- $0304d
          12366 => x"80", -- $0304e
          12367 => x"81", -- $0304f
          12368 => x"81", -- $03050
          12369 => x"80", -- $03051
          12370 => x"81", -- $03052
          12371 => x"80", -- $03053
          12372 => x"80", -- $03054
          12373 => x"81", -- $03055
          12374 => x"80", -- $03056
          12375 => x"80", -- $03057
          12376 => x"80", -- $03058
          12377 => x"80", -- $03059
          12378 => x"80", -- $0305a
          12379 => x"80", -- $0305b
          12380 => x"80", -- $0305c
          12381 => x"80", -- $0305d
          12382 => x"80", -- $0305e
          12383 => x"7f", -- $0305f
          12384 => x"80", -- $03060
          12385 => x"80", -- $03061
          12386 => x"80", -- $03062
          12387 => x"80", -- $03063
          12388 => x"80", -- $03064
          12389 => x"80", -- $03065
          12390 => x"80", -- $03066
          12391 => x"80", -- $03067
          12392 => x"80", -- $03068
          12393 => x"80", -- $03069
          12394 => x"80", -- $0306a
          12395 => x"80", -- $0306b
          12396 => x"80", -- $0306c
          12397 => x"80", -- $0306d
          12398 => x"7f", -- $0306e
          12399 => x"80", -- $0306f
          12400 => x"80", -- $03070
          12401 => x"80", -- $03071
          12402 => x"80", -- $03072
          12403 => x"80", -- $03073
          12404 => x"80", -- $03074
          12405 => x"81", -- $03075
          12406 => x"81", -- $03076
          12407 => x"80", -- $03077
          12408 => x"82", -- $03078
          12409 => x"81", -- $03079
          12410 => x"82", -- $0307a
          12411 => x"82", -- $0307b
          12412 => x"81", -- $0307c
          12413 => x"81", -- $0307d
          12414 => x"82", -- $0307e
          12415 => x"82", -- $0307f
          12416 => x"82", -- $03080
          12417 => x"82", -- $03081
          12418 => x"82", -- $03082
          12419 => x"82", -- $03083
          12420 => x"82", -- $03084
          12421 => x"81", -- $03085
          12422 => x"81", -- $03086
          12423 => x"82", -- $03087
          12424 => x"82", -- $03088
          12425 => x"81", -- $03089
          12426 => x"81", -- $0308a
          12427 => x"80", -- $0308b
          12428 => x"81", -- $0308c
          12429 => x"80", -- $0308d
          12430 => x"80", -- $0308e
          12431 => x"80", -- $0308f
          12432 => x"80", -- $03090
          12433 => x"80", -- $03091
          12434 => x"80", -- $03092
          12435 => x"80", -- $03093
          12436 => x"80", -- $03094
          12437 => x"80", -- $03095
          12438 => x"80", -- $03096
          12439 => x"80", -- $03097
          12440 => x"80", -- $03098
          12441 => x"80", -- $03099
          12442 => x"80", -- $0309a
          12443 => x"80", -- $0309b
          12444 => x"80", -- $0309c
          12445 => x"80", -- $0309d
          12446 => x"80", -- $0309e
          12447 => x"80", -- $0309f
          12448 => x"7f", -- $030a0
          12449 => x"80", -- $030a1
          12450 => x"80", -- $030a2
          12451 => x"80", -- $030a3
          12452 => x"80", -- $030a4
          12453 => x"7f", -- $030a5
          12454 => x"80", -- $030a6
          12455 => x"80", -- $030a7
          12456 => x"80", -- $030a8
          12457 => x"80", -- $030a9
          12458 => x"80", -- $030aa
          12459 => x"80", -- $030ab
          12460 => x"80", -- $030ac
          12461 => x"80", -- $030ad
          12462 => x"80", -- $030ae
          12463 => x"80", -- $030af
          12464 => x"80", -- $030b0
          12465 => x"80", -- $030b1
          12466 => x"80", -- $030b2
          12467 => x"80", -- $030b3
          12468 => x"7f", -- $030b4
          12469 => x"80", -- $030b5
          12470 => x"80", -- $030b6
          12471 => x"80", -- $030b7
          12472 => x"7f", -- $030b8
          12473 => x"80", -- $030b9
          12474 => x"7f", -- $030ba
          12475 => x"7f", -- $030bb
          12476 => x"80", -- $030bc
          12477 => x"80", -- $030bd
          12478 => x"7f", -- $030be
          12479 => x"7f", -- $030bf
          12480 => x"80", -- $030c0
          12481 => x"80", -- $030c1
          12482 => x"7f", -- $030c2
          12483 => x"7f", -- $030c3
          12484 => x"80", -- $030c4
          12485 => x"80", -- $030c5
          12486 => x"80", -- $030c6
          12487 => x"80", -- $030c7
          12488 => x"80", -- $030c8
          12489 => x"7f", -- $030c9
          12490 => x"7f", -- $030ca
          12491 => x"80", -- $030cb
          12492 => x"80", -- $030cc
          12493 => x"80", -- $030cd
          12494 => x"80", -- $030ce
          12495 => x"7f", -- $030cf
          12496 => x"7f", -- $030d0
          12497 => x"7f", -- $030d1
          12498 => x"7f", -- $030d2
          12499 => x"80", -- $030d3
          12500 => x"7f", -- $030d4
          12501 => x"7e", -- $030d5
          12502 => x"7f", -- $030d6
          12503 => x"7f", -- $030d7
          12504 => x"7f", -- $030d8
          12505 => x"7e", -- $030d9
          12506 => x"7e", -- $030da
          12507 => x"7e", -- $030db
          12508 => x"7f", -- $030dc
          12509 => x"7f", -- $030dd
          12510 => x"7e", -- $030de
          12511 => x"7e", -- $030df
          12512 => x"7e", -- $030e0
          12513 => x"7e", -- $030e1
          12514 => x"7e", -- $030e2
          12515 => x"7e", -- $030e3
          12516 => x"7e", -- $030e4
          12517 => x"7e", -- $030e5
          12518 => x"7e", -- $030e6
          12519 => x"7e", -- $030e7
          12520 => x"7e", -- $030e8
          12521 => x"7f", -- $030e9
          12522 => x"7f", -- $030ea
          12523 => x"7e", -- $030eb
          12524 => x"7e", -- $030ec
          12525 => x"7f", -- $030ed
          12526 => x"7f", -- $030ee
          12527 => x"7f", -- $030ef
          12528 => x"80", -- $030f0
          12529 => x"80", -- $030f1
          12530 => x"80", -- $030f2
          12531 => x"80", -- $030f3
          12532 => x"80", -- $030f4
          12533 => x"80", -- $030f5
          12534 => x"80", -- $030f6
          12535 => x"80", -- $030f7
          12536 => x"80", -- $030f8
          12537 => x"7f", -- $030f9
          12538 => x"7f", -- $030fa
          12539 => x"7f", -- $030fb
          12540 => x"7f", -- $030fc
          12541 => x"7f", -- $030fd
          12542 => x"7f", -- $030fe
          12543 => x"7f", -- $030ff
          12544 => x"7f", -- $03100
          12545 => x"7f", -- $03101
          12546 => x"7f", -- $03102
          12547 => x"7f", -- $03103
          12548 => x"80", -- $03104
          12549 => x"7f", -- $03105
          12550 => x"7f", -- $03106
          12551 => x"7f", -- $03107
          12552 => x"7f", -- $03108
          12553 => x"7f", -- $03109
          12554 => x"7f", -- $0310a
          12555 => x"7f", -- $0310b
          12556 => x"7f", -- $0310c
          12557 => x"7f", -- $0310d
          12558 => x"7f", -- $0310e
          12559 => x"7f", -- $0310f
          12560 => x"7f", -- $03110
          12561 => x"7f", -- $03111
          12562 => x"7f", -- $03112
          12563 => x"7f", -- $03113
          12564 => x"7f", -- $03114
          12565 => x"7f", -- $03115
          12566 => x"7f", -- $03116
          12567 => x"7f", -- $03117
          12568 => x"7f", -- $03118
          12569 => x"7f", -- $03119
          12570 => x"7f", -- $0311a
          12571 => x"7f", -- $0311b
          12572 => x"7f", -- $0311c
          12573 => x"7f", -- $0311d
          12574 => x"7f", -- $0311e
          12575 => x"7f", -- $0311f
          12576 => x"7f", -- $03120
          12577 => x"7f", -- $03121
          12578 => x"7f", -- $03122
          12579 => x"7f", -- $03123
          12580 => x"7f", -- $03124
          12581 => x"7f", -- $03125
          12582 => x"80", -- $03126
          12583 => x"80", -- $03127
          12584 => x"80", -- $03128
          12585 => x"80", -- $03129
          12586 => x"80", -- $0312a
          12587 => x"80", -- $0312b
          12588 => x"80", -- $0312c
          12589 => x"80", -- $0312d
          12590 => x"80", -- $0312e
          12591 => x"80", -- $0312f
          12592 => x"80", -- $03130
          12593 => x"80", -- $03131
          12594 => x"80", -- $03132
          12595 => x"80", -- $03133
          12596 => x"80", -- $03134
          12597 => x"80", -- $03135
          12598 => x"80", -- $03136
          12599 => x"80", -- $03137
          12600 => x"80", -- $03138
          12601 => x"80", -- $03139
          12602 => x"80", -- $0313a
          12603 => x"80", -- $0313b
          12604 => x"80", -- $0313c
          12605 => x"80", -- $0313d
          12606 => x"80", -- $0313e
          12607 => x"80", -- $0313f
          12608 => x"80", -- $03140
          12609 => x"80", -- $03141
          12610 => x"80", -- $03142
          12611 => x"80", -- $03143
          12612 => x"80", -- $03144
          12613 => x"80", -- $03145
          12614 => x"80", -- $03146
          12615 => x"80", -- $03147
          12616 => x"80", -- $03148
          12617 => x"80", -- $03149
          12618 => x"80", -- $0314a
          12619 => x"80", -- $0314b
          12620 => x"80", -- $0314c
          12621 => x"80", -- $0314d
          12622 => x"80", -- $0314e
          12623 => x"7f", -- $0314f
          12624 => x"7f", -- $03150
          12625 => x"7f", -- $03151
          12626 => x"7f", -- $03152
          12627 => x"7f", -- $03153
          12628 => x"7f", -- $03154
          12629 => x"7f", -- $03155
          12630 => x"7f", -- $03156
          12631 => x"7f", -- $03157
          12632 => x"7f", -- $03158
          12633 => x"7f", -- $03159
          12634 => x"7f", -- $0315a
          12635 => x"7f", -- $0315b
          12636 => x"7f", -- $0315c
          12637 => x"80", -- $0315d
          12638 => x"80", -- $0315e
          12639 => x"80", -- $0315f
          12640 => x"80", -- $03160
          12641 => x"80", -- $03161
          12642 => x"80", -- $03162
          12643 => x"80", -- $03163
          12644 => x"80", -- $03164
          12645 => x"80", -- $03165
          12646 => x"80", -- $03166
          12647 => x"80", -- $03167
          12648 => x"80", -- $03168
          12649 => x"80", -- $03169
          12650 => x"80", -- $0316a
          12651 => x"80", -- $0316b
          12652 => x"80", -- $0316c
          12653 => x"80", -- $0316d
          12654 => x"80", -- $0316e
          12655 => x"80", -- $0316f
          12656 => x"80", -- $03170
          12657 => x"80", -- $03171
          12658 => x"80", -- $03172
          12659 => x"80", -- $03173
          12660 => x"80", -- $03174
          12661 => x"80", -- $03175
          12662 => x"80", -- $03176
          12663 => x"80", -- $03177
          12664 => x"7f", -- $03178
          12665 => x"7f", -- $03179
          12666 => x"7f", -- $0317a
          12667 => x"7f", -- $0317b
          12668 => x"7f", -- $0317c
          12669 => x"7f", -- $0317d
          12670 => x"7f", -- $0317e
          12671 => x"7f", -- $0317f
          12672 => x"7f", -- $03180
          12673 => x"7f", -- $03181
          12674 => x"7f", -- $03182
          12675 => x"7f", -- $03183
          12676 => x"80", -- $03184
          12677 => x"80", -- $03185
          12678 => x"80", -- $03186
          12679 => x"80", -- $03187
          12680 => x"80", -- $03188
          12681 => x"80", -- $03189
          12682 => x"80", -- $0318a
          12683 => x"80", -- $0318b
          12684 => x"80", -- $0318c
          12685 => x"80", -- $0318d
          12686 => x"80", -- $0318e
          12687 => x"80", -- $0318f
          12688 => x"80", -- $03190
          12689 => x"80", -- $03191
          12690 => x"7f", -- $03192
          12691 => x"7f", -- $03193
          12692 => x"7e", -- $03194
          12693 => x"7e", -- $03195
          12694 => x"7e", -- $03196
          12695 => x"7e", -- $03197
          12696 => x"7e", -- $03198
          12697 => x"7e", -- $03199
          12698 => x"7e", -- $0319a
          12699 => x"7e", -- $0319b
          12700 => x"7f", -- $0319c
          12701 => x"7f", -- $0319d
          12702 => x"7f", -- $0319e
          12703 => x"80", -- $0319f
          12704 => x"80", -- $031a0
          12705 => x"7f", -- $031a1
          12706 => x"7f", -- $031a2
          12707 => x"7f", -- $031a3
          12708 => x"7f", -- $031a4
          12709 => x"80", -- $031a5
          12710 => x"80", -- $031a6
          12711 => x"80", -- $031a7
          12712 => x"80", -- $031a8
          12713 => x"80", -- $031a9
          12714 => x"80", -- $031aa
          12715 => x"80", -- $031ab
          12716 => x"80", -- $031ac
          12717 => x"80", -- $031ad
          12718 => x"80", -- $031ae
          12719 => x"80", -- $031af
          12720 => x"80", -- $031b0
          12721 => x"80", -- $031b1
          12722 => x"80", -- $031b2
          12723 => x"7f", -- $031b3
          12724 => x"80", -- $031b4
          12725 => x"80", -- $031b5
          12726 => x"80", -- $031b6
          12727 => x"80", -- $031b7
          12728 => x"7f", -- $031b8
          12729 => x"80", -- $031b9
          12730 => x"80", -- $031ba
          12731 => x"7f", -- $031bb
          12732 => x"7f", -- $031bc
          12733 => x"7f", -- $031bd
          12734 => x"7f", -- $031be
          12735 => x"7f", -- $031bf
          12736 => x"7f", -- $031c0
          12737 => x"7f", -- $031c1
          12738 => x"80", -- $031c2
          12739 => x"80", -- $031c3
          12740 => x"80", -- $031c4
          12741 => x"80", -- $031c5
          12742 => x"80", -- $031c6
          12743 => x"80", -- $031c7
          12744 => x"80", -- $031c8
          12745 => x"80", -- $031c9
          12746 => x"80", -- $031ca
          12747 => x"80", -- $031cb
          12748 => x"80", -- $031cc
          12749 => x"7f", -- $031cd
          12750 => x"7f", -- $031ce
          12751 => x"7f", -- $031cf
          12752 => x"7f", -- $031d0
          12753 => x"80", -- $031d1
          12754 => x"80", -- $031d2
          12755 => x"80", -- $031d3
          12756 => x"80", -- $031d4
          12757 => x"80", -- $031d5
          12758 => x"7f", -- $031d6
          12759 => x"7f", -- $031d7
          12760 => x"80", -- $031d8
          12761 => x"80", -- $031d9
          12762 => x"80", -- $031da
          12763 => x"80", -- $031db
          12764 => x"80", -- $031dc
          12765 => x"80", -- $031dd
          12766 => x"80", -- $031de
          12767 => x"80", -- $031df
          12768 => x"80", -- $031e0
          12769 => x"80", -- $031e1
          12770 => x"80", -- $031e2
          12771 => x"80", -- $031e3
          12772 => x"80", -- $031e4
          12773 => x"80", -- $031e5
          12774 => x"80", -- $031e6
          12775 => x"80", -- $031e7
          12776 => x"80", -- $031e8
          12777 => x"80", -- $031e9
          12778 => x"80", -- $031ea
          12779 => x"80", -- $031eb
          12780 => x"80", -- $031ec
          12781 => x"80", -- $031ed
          12782 => x"80", -- $031ee
          12783 => x"80", -- $031ef
          12784 => x"80", -- $031f0
          12785 => x"80", -- $031f1
          12786 => x"80", -- $031f2
          12787 => x"80", -- $031f3
          12788 => x"7f", -- $031f4
          12789 => x"7f", -- $031f5
          12790 => x"7f", -- $031f6
          12791 => x"7f", -- $031f7
          12792 => x"7f", -- $031f8
          12793 => x"7f", -- $031f9
          12794 => x"80", -- $031fa
          12795 => x"80", -- $031fb
          12796 => x"80", -- $031fc
          12797 => x"80", -- $031fd
          12798 => x"80", -- $031fe
          12799 => x"80", -- $031ff
          12800 => x"80", -- $03200
          12801 => x"80", -- $03201
          12802 => x"80", -- $03202
          12803 => x"80", -- $03203
          12804 => x"80", -- $03204
          12805 => x"80", -- $03205
          12806 => x"80", -- $03206
          12807 => x"80", -- $03207
          12808 => x"80", -- $03208
          12809 => x"80", -- $03209
          12810 => x"80", -- $0320a
          12811 => x"80", -- $0320b
          12812 => x"80", -- $0320c
          12813 => x"80", -- $0320d
          12814 => x"80", -- $0320e
          12815 => x"80", -- $0320f
          12816 => x"80", -- $03210
          12817 => x"80", -- $03211
          12818 => x"80", -- $03212
          12819 => x"80", -- $03213
          12820 => x"80", -- $03214
          12821 => x"80", -- $03215
          12822 => x"80", -- $03216
          12823 => x"80", -- $03217
          12824 => x"80", -- $03218
          12825 => x"80", -- $03219
          12826 => x"80", -- $0321a
          12827 => x"80", -- $0321b
          12828 => x"80", -- $0321c
          12829 => x"80", -- $0321d
          12830 => x"80", -- $0321e
          12831 => x"80", -- $0321f
          12832 => x"80", -- $03220
          12833 => x"80", -- $03221
          12834 => x"80", -- $03222
          12835 => x"80", -- $03223
          12836 => x"80", -- $03224
          12837 => x"80", -- $03225
          12838 => x"80", -- $03226
          12839 => x"80", -- $03227
          12840 => x"80", -- $03228
          12841 => x"80", -- $03229
          12842 => x"80", -- $0322a
          12843 => x"80", -- $0322b
          12844 => x"80", -- $0322c
          12845 => x"80", -- $0322d
          12846 => x"80", -- $0322e
          12847 => x"81", -- $0322f
          12848 => x"81", -- $03230
          12849 => x"81", -- $03231
          12850 => x"81", -- $03232
          12851 => x"81", -- $03233
          12852 => x"81", -- $03234
          12853 => x"81", -- $03235
          12854 => x"81", -- $03236
          12855 => x"80", -- $03237
          12856 => x"80", -- $03238
          12857 => x"80", -- $03239
          12858 => x"80", -- $0323a
          12859 => x"80", -- $0323b
          12860 => x"80", -- $0323c
          12861 => x"80", -- $0323d
          12862 => x"80", -- $0323e
          12863 => x"80", -- $0323f
          12864 => x"80", -- $03240
          12865 => x"80", -- $03241
          12866 => x"81", -- $03242
          12867 => x"81", -- $03243
          12868 => x"82", -- $03244
          12869 => x"82", -- $03245
          12870 => x"82", -- $03246
          12871 => x"82", -- $03247
          12872 => x"82", -- $03248
          12873 => x"81", -- $03249
          12874 => x"81", -- $0324a
          12875 => x"81", -- $0324b
          12876 => x"81", -- $0324c
          12877 => x"81", -- $0324d
          12878 => x"81", -- $0324e
          12879 => x"81", -- $0324f
          12880 => x"80", -- $03250
          12881 => x"80", -- $03251
          12882 => x"81", -- $03252
          12883 => x"81", -- $03253
          12884 => x"81", -- $03254
          12885 => x"81", -- $03255
          12886 => x"81", -- $03256
          12887 => x"81", -- $03257
          12888 => x"81", -- $03258
          12889 => x"80", -- $03259
          12890 => x"80", -- $0325a
          12891 => x"80", -- $0325b
          12892 => x"80", -- $0325c
          12893 => x"80", -- $0325d
          12894 => x"80", -- $0325e
          12895 => x"80", -- $0325f
          12896 => x"80", -- $03260
          12897 => x"81", -- $03261
          12898 => x"81", -- $03262
          12899 => x"81", -- $03263
          12900 => x"81", -- $03264
          12901 => x"81", -- $03265
          12902 => x"81", -- $03266
          12903 => x"81", -- $03267
          12904 => x"80", -- $03268
          12905 => x"80", -- $03269
          12906 => x"80", -- $0326a
          12907 => x"81", -- $0326b
          12908 => x"81", -- $0326c
          12909 => x"81", -- $0326d
          12910 => x"81", -- $0326e
          12911 => x"81", -- $0326f
          12912 => x"80", -- $03270
          12913 => x"80", -- $03271
          12914 => x"81", -- $03272
          12915 => x"81", -- $03273
          12916 => x"81", -- $03274
          12917 => x"81", -- $03275
          12918 => x"81", -- $03276
          12919 => x"81", -- $03277
          12920 => x"81", -- $03278
          12921 => x"81", -- $03279
          12922 => x"81", -- $0327a
          12923 => x"81", -- $0327b
          12924 => x"81", -- $0327c
          12925 => x"81", -- $0327d
          12926 => x"81", -- $0327e
          12927 => x"80", -- $0327f
          12928 => x"80", -- $03280
          12929 => x"80", -- $03281
          12930 => x"80", -- $03282
          12931 => x"80", -- $03283
          12932 => x"80", -- $03284
          12933 => x"80", -- $03285
          12934 => x"80", -- $03286
          12935 => x"80", -- $03287
          12936 => x"80", -- $03288
          12937 => x"80", -- $03289
          12938 => x"80", -- $0328a
          12939 => x"80", -- $0328b
          12940 => x"80", -- $0328c
          12941 => x"80", -- $0328d
          12942 => x"80", -- $0328e
          12943 => x"80", -- $0328f
          12944 => x"80", -- $03290
          12945 => x"80", -- $03291
          12946 => x"80", -- $03292
          12947 => x"80", -- $03293
          12948 => x"80", -- $03294
          12949 => x"80", -- $03295
          12950 => x"80", -- $03296
          12951 => x"80", -- $03297
          12952 => x"80", -- $03298
          12953 => x"80", -- $03299
          12954 => x"80", -- $0329a
          12955 => x"80", -- $0329b
          12956 => x"80", -- $0329c
          12957 => x"80", -- $0329d
          12958 => x"80", -- $0329e
          12959 => x"80", -- $0329f
          12960 => x"80", -- $032a0
          12961 => x"80", -- $032a1
          12962 => x"80", -- $032a2
          12963 => x"80", -- $032a3
          12964 => x"80", -- $032a4
          12965 => x"80", -- $032a5
          12966 => x"80", -- $032a6
          12967 => x"80", -- $032a7
          12968 => x"80", -- $032a8
          12969 => x"80", -- $032a9
          12970 => x"81", -- $032aa
          12971 => x"81", -- $032ab
          12972 => x"81", -- $032ac
          12973 => x"81", -- $032ad
          12974 => x"81", -- $032ae
          12975 => x"81", -- $032af
          12976 => x"80", -- $032b0
          12977 => x"80", -- $032b1
          12978 => x"80", -- $032b2
          12979 => x"80", -- $032b3
          12980 => x"80", -- $032b4
          12981 => x"80", -- $032b5
          12982 => x"80", -- $032b6
          12983 => x"80", -- $032b7
          12984 => x"80", -- $032b8
          12985 => x"80", -- $032b9
          12986 => x"80", -- $032ba
          12987 => x"80", -- $032bb
          12988 => x"80", -- $032bc
          12989 => x"80", -- $032bd
          12990 => x"80", -- $032be
          12991 => x"80", -- $032bf
          12992 => x"80", -- $032c0
          12993 => x"80", -- $032c1
          12994 => x"80", -- $032c2
          12995 => x"80", -- $032c3
          12996 => x"80", -- $032c4
          12997 => x"80", -- $032c5
          12998 => x"80", -- $032c6
          12999 => x"80", -- $032c7
          13000 => x"80", -- $032c8
          13001 => x"80", -- $032c9
          13002 => x"81", -- $032ca
          13003 => x"81", -- $032cb
          13004 => x"81", -- $032cc
          13005 => x"81", -- $032cd
          13006 => x"81", -- $032ce
          13007 => x"82", -- $032cf
          13008 => x"82", -- $032d0
          13009 => x"83", -- $032d1
          13010 => x"83", -- $032d2
          13011 => x"84", -- $032d3
          13012 => x"84", -- $032d4
          13013 => x"84", -- $032d5
          13014 => x"85", -- $032d6
          13015 => x"85", -- $032d7
          13016 => x"84", -- $032d8
          13017 => x"84", -- $032d9
          13018 => x"84", -- $032da
          13019 => x"83", -- $032db
          13020 => x"83", -- $032dc
          13021 => x"82", -- $032dd
          13022 => x"82", -- $032de
          13023 => x"81", -- $032df
          13024 => x"81", -- $032e0
          13025 => x"80", -- $032e1
          13026 => x"80", -- $032e2
          13027 => x"7f", -- $032e3
          13028 => x"7f", -- $032e4
          13029 => x"7e", -- $032e5
          13030 => x"7e", -- $032e6
          13031 => x"7d", -- $032e7
          13032 => x"7d", -- $032e8
          13033 => x"7d", -- $032e9
          13034 => x"7e", -- $032ea
          13035 => x"7e", -- $032eb
          13036 => x"7e", -- $032ec
          13037 => x"7f", -- $032ed
          13038 => x"7f", -- $032ee
          13039 => x"80", -- $032ef
          13040 => x"80", -- $032f0
          13041 => x"80", -- $032f1
          13042 => x"80", -- $032f2
          13043 => x"80", -- $032f3
          13044 => x"81", -- $032f4
          13045 => x"81", -- $032f5
          13046 => x"81", -- $032f6
          13047 => x"82", -- $032f7
          13048 => x"82", -- $032f8
          13049 => x"82", -- $032f9
          13050 => x"82", -- $032fa
          13051 => x"82", -- $032fb
          13052 => x"82", -- $032fc
          13053 => x"82", -- $032fd
          13054 => x"82", -- $032fe
          13055 => x"82", -- $032ff
          13056 => x"83", -- $03300
          13057 => x"84", -- $03301
          13058 => x"84", -- $03302
          13059 => x"85", -- $03303
          13060 => x"85", -- $03304
          13061 => x"86", -- $03305
          13062 => x"86", -- $03306
          13063 => x"86", -- $03307
          13064 => x"86", -- $03308
          13065 => x"85", -- $03309
          13066 => x"85", -- $0330a
          13067 => x"84", -- $0330b
          13068 => x"84", -- $0330c
          13069 => x"83", -- $0330d
          13070 => x"82", -- $0330e
          13071 => x"81", -- $0330f
          13072 => x"81", -- $03310
          13073 => x"80", -- $03311
          13074 => x"80", -- $03312
          13075 => x"7f", -- $03313
          13076 => x"7e", -- $03314
          13077 => x"7d", -- $03315
          13078 => x"7c", -- $03316
          13079 => x"7b", -- $03317
          13080 => x"7b", -- $03318
          13081 => x"7b", -- $03319
          13082 => x"7b", -- $0331a
          13083 => x"7c", -- $0331b
          13084 => x"7d", -- $0331c
          13085 => x"7e", -- $0331d
          13086 => x"7f", -- $0331e
          13087 => x"80", -- $0331f
          13088 => x"80", -- $03320
          13089 => x"81", -- $03321
          13090 => x"81", -- $03322
          13091 => x"82", -- $03323
          13092 => x"82", -- $03324
          13093 => x"83", -- $03325
          13094 => x"83", -- $03326
          13095 => x"83", -- $03327
          13096 => x"82", -- $03328
          13097 => x"81", -- $03329
          13098 => x"80", -- $0332a
          13099 => x"7f", -- $0332b
          13100 => x"7e", -- $0332c
          13101 => x"7c", -- $0332d
          13102 => x"7b", -- $0332e
          13103 => x"7b", -- $0332f
          13104 => x"7b", -- $03330
          13105 => x"7c", -- $03331
          13106 => x"7c", -- $03332
          13107 => x"7e", -- $03333
          13108 => x"7f", -- $03334
          13109 => x"80", -- $03335
          13110 => x"80", -- $03336
          13111 => x"82", -- $03337
          13112 => x"83", -- $03338
          13113 => x"83", -- $03339
          13114 => x"83", -- $0333a
          13115 => x"84", -- $0333b
          13116 => x"84", -- $0333c
          13117 => x"83", -- $0333d
          13118 => x"83", -- $0333e
          13119 => x"83", -- $0333f
          13120 => x"83", -- $03340
          13121 => x"83", -- $03341
          13122 => x"84", -- $03342
          13123 => x"84", -- $03343
          13124 => x"84", -- $03344
          13125 => x"83", -- $03345
          13126 => x"83", -- $03346
          13127 => x"82", -- $03347
          13128 => x"82", -- $03348
          13129 => x"82", -- $03349
          13130 => x"82", -- $0334a
          13131 => x"82", -- $0334b
          13132 => x"83", -- $0334c
          13133 => x"83", -- $0334d
          13134 => x"83", -- $0334e
          13135 => x"82", -- $0334f
          13136 => x"80", -- $03350
          13137 => x"7f", -- $03351
          13138 => x"7d", -- $03352
          13139 => x"7b", -- $03353
          13140 => x"7a", -- $03354
          13141 => x"79", -- $03355
          13142 => x"79", -- $03356
          13143 => x"79", -- $03357
          13144 => x"7a", -- $03358
          13145 => x"7b", -- $03359
          13146 => x"7d", -- $0335a
          13147 => x"7e", -- $0335b
          13148 => x"7e", -- $0335c
          13149 => x"7f", -- $0335d
          13150 => x"7f", -- $0335e
          13151 => x"80", -- $0335f
          13152 => x"80", -- $03360
          13153 => x"80", -- $03361
          13154 => x"81", -- $03362
          13155 => x"81", -- $03363
          13156 => x"81", -- $03364
          13157 => x"80", -- $03365
          13158 => x"80", -- $03366
          13159 => x"7e", -- $03367
          13160 => x"7d", -- $03368
          13161 => x"7c", -- $03369
          13162 => x"7c", -- $0336a
          13163 => x"7c", -- $0336b
          13164 => x"7c", -- $0336c
          13165 => x"7d", -- $0336d
          13166 => x"7f", -- $0336e
          13167 => x"80", -- $0336f
          13168 => x"81", -- $03370
          13169 => x"83", -- $03371
          13170 => x"85", -- $03372
          13171 => x"87", -- $03373
          13172 => x"88", -- $03374
          13173 => x"8a", -- $03375
          13174 => x"8b", -- $03376
          13175 => x"8b", -- $03377
          13176 => x"8b", -- $03378
          13177 => x"89", -- $03379
          13178 => x"86", -- $0337a
          13179 => x"84", -- $0337b
          13180 => x"82", -- $0337c
          13181 => x"81", -- $0337d
          13182 => x"81", -- $0337e
          13183 => x"80", -- $0337f
          13184 => x"80", -- $03380
          13185 => x"80", -- $03381
          13186 => x"7f", -- $03382
          13187 => x"7d", -- $03383
          13188 => x"7a", -- $03384
          13189 => x"78", -- $03385
          13190 => x"76", -- $03386
          13191 => x"75", -- $03387
          13192 => x"75", -- $03388
          13193 => x"77", -- $03389
          13194 => x"79", -- $0338a
          13195 => x"7b", -- $0338b
          13196 => x"7e", -- $0338c
          13197 => x"80", -- $0338d
          13198 => x"81", -- $0338e
          13199 => x"82", -- $0338f
          13200 => x"83", -- $03390
          13201 => x"83", -- $03391
          13202 => x"84", -- $03392
          13203 => x"85", -- $03393
          13204 => x"86", -- $03394
          13205 => x"87", -- $03395
          13206 => x"86", -- $03396
          13207 => x"84", -- $03397
          13208 => x"81", -- $03398
          13209 => x"7f", -- $03399
          13210 => x"7b", -- $0339a
          13211 => x"78", -- $0339b
          13212 => x"76", -- $0339c
          13213 => x"75", -- $0339d
          13214 => x"75", -- $0339e
          13215 => x"76", -- $0339f
          13216 => x"77", -- $033a0
          13217 => x"79", -- $033a1
          13218 => x"7a", -- $033a2
          13219 => x"7c", -- $033a3
          13220 => x"7e", -- $033a4
          13221 => x"80", -- $033a5
          13222 => x"82", -- $033a6
          13223 => x"84", -- $033a7
          13224 => x"85", -- $033a8
          13225 => x"85", -- $033a9
          13226 => x"85", -- $033aa
          13227 => x"84", -- $033ab
          13228 => x"83", -- $033ac
          13229 => x"81", -- $033ad
          13230 => x"80", -- $033ae
          13231 => x"80", -- $033af
          13232 => x"80", -- $033b0
          13233 => x"80", -- $033b1
          13234 => x"81", -- $033b2
          13235 => x"83", -- $033b3
          13236 => x"83", -- $033b4
          13237 => x"82", -- $033b5
          13238 => x"81", -- $033b6
          13239 => x"80", -- $033b7
          13240 => x"80", -- $033b8
          13241 => x"80", -- $033b9
          13242 => x"81", -- $033ba
          13243 => x"83", -- $033bb
          13244 => x"85", -- $033bc
          13245 => x"85", -- $033bd
          13246 => x"84", -- $033be
          13247 => x"82", -- $033bf
          13248 => x"80", -- $033c0
          13249 => x"7d", -- $033c1
          13250 => x"7b", -- $033c2
          13251 => x"7a", -- $033c3
          13252 => x"7a", -- $033c4
          13253 => x"7b", -- $033c5
          13254 => x"7d", -- $033c6
          13255 => x"7d", -- $033c7
          13256 => x"7d", -- $033c8
          13257 => x"7d", -- $033c9
          13258 => x"7d", -- $033ca
          13259 => x"7d", -- $033cb
          13260 => x"7e", -- $033cc
          13261 => x"80", -- $033cd
          13262 => x"81", -- $033ce
          13263 => x"83", -- $033cf
          13264 => x"85", -- $033d0
          13265 => x"84", -- $033d1
          13266 => x"83", -- $033d2
          13267 => x"81", -- $033d3
          13268 => x"7f", -- $033d4
          13269 => x"7c", -- $033d5
          13270 => x"7a", -- $033d6
          13271 => x"79", -- $033d7
          13272 => x"79", -- $033d8
          13273 => x"78", -- $033d9
          13274 => x"78", -- $033da
          13275 => x"77", -- $033db
          13276 => x"76", -- $033dc
          13277 => x"76", -- $033dd
          13278 => x"76", -- $033de
          13279 => x"79", -- $033df
          13280 => x"7c", -- $033e0
          13281 => x"80", -- $033e1
          13282 => x"83", -- $033e2
          13283 => x"85", -- $033e3
          13284 => x"87", -- $033e4
          13285 => x"88", -- $033e5
          13286 => x"88", -- $033e6
          13287 => x"88", -- $033e7
          13288 => x"88", -- $033e8
          13289 => x"88", -- $033e9
          13290 => x"89", -- $033ea
          13291 => x"89", -- $033eb
          13292 => x"87", -- $033ec
          13293 => x"83", -- $033ed
          13294 => x"80", -- $033ee
          13295 => x"7c", -- $033ef
          13296 => x"79", -- $033f0
          13297 => x"79", -- $033f1
          13298 => x"7c", -- $033f2
          13299 => x"7f", -- $033f3
          13300 => x"81", -- $033f4
          13301 => x"82", -- $033f5
          13302 => x"81", -- $033f6
          13303 => x"80", -- $033f7
          13304 => x"7e", -- $033f8
          13305 => x"7c", -- $033f9
          13306 => x"7d", -- $033fa
          13307 => x"7e", -- $033fb
          13308 => x"80", -- $033fc
          13309 => x"80", -- $033fd
          13310 => x"80", -- $033fe
          13311 => x"7f", -- $033ff
          13312 => x"7d", -- $03400
          13313 => x"7c", -- $03401
          13314 => x"7c", -- $03402
          13315 => x"7d", -- $03403
          13316 => x"7f", -- $03404
          13317 => x"80", -- $03405
          13318 => x"82", -- $03406
          13319 => x"82", -- $03407
          13320 => x"82", -- $03408
          13321 => x"81", -- $03409
          13322 => x"80", -- $0340a
          13323 => x"80", -- $0340b
          13324 => x"7f", -- $0340c
          13325 => x"80", -- $0340d
          13326 => x"7f", -- $0340e
          13327 => x"7e", -- $0340f
          13328 => x"7c", -- $03410
          13329 => x"7a", -- $03411
          13330 => x"78", -- $03412
          13331 => x"78", -- $03413
          13332 => x"79", -- $03414
          13333 => x"7b", -- $03415
          13334 => x"7d", -- $03416
          13335 => x"7f", -- $03417
          13336 => x"80", -- $03418
          13337 => x"80", -- $03419
          13338 => x"80", -- $0341a
          13339 => x"81", -- $0341b
          13340 => x"81", -- $0341c
          13341 => x"82", -- $0341d
          13342 => x"82", -- $0341e
          13343 => x"82", -- $0341f
          13344 => x"80", -- $03420
          13345 => x"7f", -- $03421
          13346 => x"7d", -- $03422
          13347 => x"7d", -- $03423
          13348 => x"7d", -- $03424
          13349 => x"7f", -- $03425
          13350 => x"80", -- $03426
          13351 => x"82", -- $03427
          13352 => x"82", -- $03428
          13353 => x"81", -- $03429
          13354 => x"80", -- $0342a
          13355 => x"80", -- $0342b
          13356 => x"81", -- $0342c
          13357 => x"83", -- $0342d
          13358 => x"85", -- $0342e
          13359 => x"86", -- $0342f
          13360 => x"86", -- $03430
          13361 => x"84", -- $03431
          13362 => x"81", -- $03432
          13363 => x"80", -- $03433
          13364 => x"7e", -- $03434
          13365 => x"7d", -- $03435
          13366 => x"7d", -- $03436
          13367 => x"7e", -- $03437
          13368 => x"7e", -- $03438
          13369 => x"7c", -- $03439
          13370 => x"7b", -- $0343a
          13371 => x"7a", -- $0343b
          13372 => x"7a", -- $0343c
          13373 => x"7b", -- $0343d
          13374 => x"7e", -- $0343e
          13375 => x"80", -- $0343f
          13376 => x"80", -- $03440
          13377 => x"81", -- $03441
          13378 => x"80", -- $03442
          13379 => x"80", -- $03443
          13380 => x"7f", -- $03444
          13381 => x"7e", -- $03445
          13382 => x"7f", -- $03446
          13383 => x"7e", -- $03447
          13384 => x"7d", -- $03448
          13385 => x"7b", -- $03449
          13386 => x"79", -- $0344a
          13387 => x"77", -- $0344b
          13388 => x"77", -- $0344c
          13389 => x"77", -- $0344d
          13390 => x"78", -- $0344e
          13391 => x"7a", -- $0344f
          13392 => x"7b", -- $03450
          13393 => x"7b", -- $03451
          13394 => x"7c", -- $03452
          13395 => x"7d", -- $03453
          13396 => x"80", -- $03454
          13397 => x"81", -- $03455
          13398 => x"84", -- $03456
          13399 => x"86", -- $03457
          13400 => x"86", -- $03458
          13401 => x"86", -- $03459
          13402 => x"86", -- $0345a
          13403 => x"86", -- $0345b
          13404 => x"85", -- $0345c
          13405 => x"83", -- $0345d
          13406 => x"82", -- $0345e
          13407 => x"80", -- $0345f
          13408 => x"7f", -- $03460
          13409 => x"80", -- $03461
          13410 => x"7f", -- $03462
          13411 => x"80", -- $03463
          13412 => x"80", -- $03464
          13413 => x"80", -- $03465
          13414 => x"80", -- $03466
          13415 => x"7f", -- $03467
          13416 => x"7f", -- $03468
          13417 => x"7e", -- $03469
          13418 => x"7e", -- $0346a
          13419 => x"7d", -- $0346b
          13420 => x"7c", -- $0346c
          13421 => x"7c", -- $0346d
          13422 => x"7b", -- $0346e
          13423 => x"7b", -- $0346f
          13424 => x"7c", -- $03470
          13425 => x"7d", -- $03471
          13426 => x"7e", -- $03472
          13427 => x"80", -- $03473
          13428 => x"80", -- $03474
          13429 => x"80", -- $03475
          13430 => x"80", -- $03476
          13431 => x"81", -- $03477
          13432 => x"82", -- $03478
          13433 => x"83", -- $03479
          13434 => x"83", -- $0347a
          13435 => x"82", -- $0347b
          13436 => x"80", -- $0347c
          13437 => x"7f", -- $0347d
          13438 => x"7c", -- $0347e
          13439 => x"7b", -- $0347f
          13440 => x"7a", -- $03480
          13441 => x"7a", -- $03481
          13442 => x"7a", -- $03482
          13443 => x"7a", -- $03483
          13444 => x"7b", -- $03484
          13445 => x"7c", -- $03485
          13446 => x"7e", -- $03486
          13447 => x"80", -- $03487
          13448 => x"82", -- $03488
          13449 => x"84", -- $03489
          13450 => x"84", -- $0348a
          13451 => x"83", -- $0348b
          13452 => x"82", -- $0348c
          13453 => x"81", -- $0348d
          13454 => x"80", -- $0348e
          13455 => x"80", -- $0348f
          13456 => x"7e", -- $03490
          13457 => x"7c", -- $03491
          13458 => x"7b", -- $03492
          13459 => x"7a", -- $03493
          13460 => x"7a", -- $03494
          13461 => x"7b", -- $03495
          13462 => x"7d", -- $03496
          13463 => x"80", -- $03497
          13464 => x"82", -- $03498
          13465 => x"84", -- $03499
          13466 => x"84", -- $0349a
          13467 => x"84", -- $0349b
          13468 => x"83", -- $0349c
          13469 => x"83", -- $0349d
          13470 => x"84", -- $0349e
          13471 => x"84", -- $0349f
          13472 => x"85", -- $034a0
          13473 => x"84", -- $034a1
          13474 => x"81", -- $034a2
          13475 => x"80", -- $034a3
          13476 => x"7f", -- $034a4
          13477 => x"7d", -- $034a5
          13478 => x"7d", -- $034a6
          13479 => x"7e", -- $034a7
          13480 => x"7d", -- $034a8
          13481 => x"7d", -- $034a9
          13482 => x"7b", -- $034aa
          13483 => x"7b", -- $034ab
          13484 => x"7b", -- $034ac
          13485 => x"7d", -- $034ad
          13486 => x"80", -- $034ae
          13487 => x"81", -- $034af
          13488 => x"82", -- $034b0
          13489 => x"82", -- $034b1
          13490 => x"81", -- $034b2
          13491 => x"80", -- $034b3
          13492 => x"81", -- $034b4
          13493 => x"81", -- $034b5
          13494 => x"82", -- $034b6
          13495 => x"81", -- $034b7
          13496 => x"80", -- $034b8
          13497 => x"7d", -- $034b9
          13498 => x"7b", -- $034ba
          13499 => x"7b", -- $034bb
          13500 => x"7a", -- $034bc
          13501 => x"7a", -- $034bd
          13502 => x"7b", -- $034be
          13503 => x"7b", -- $034bf
          13504 => x"7a", -- $034c0
          13505 => x"7b", -- $034c1
          13506 => x"7c", -- $034c2
          13507 => x"7e", -- $034c3
          13508 => x"80", -- $034c4
          13509 => x"83", -- $034c5
          13510 => x"85", -- $034c6
          13511 => x"85", -- $034c7
          13512 => x"86", -- $034c8
          13513 => x"87", -- $034c9
          13514 => x"88", -- $034ca
          13515 => x"89", -- $034cb
          13516 => x"8a", -- $034cc
          13517 => x"88", -- $034cd
          13518 => x"83", -- $034ce
          13519 => x"80", -- $034cf
          13520 => x"7e", -- $034d0
          13521 => x"7c", -- $034d1
          13522 => x"7e", -- $034d2
          13523 => x"7f", -- $034d3
          13524 => x"80", -- $034d4
          13525 => x"7f", -- $034d5
          13526 => x"7d", -- $034d6
          13527 => x"7e", -- $034d7
          13528 => x"7e", -- $034d8
          13529 => x"7f", -- $034d9
          13530 => x"80", -- $034da
          13531 => x"80", -- $034db
          13532 => x"7f", -- $034dc
          13533 => x"7d", -- $034dd
          13534 => x"7c", -- $034de
          13535 => x"7c", -- $034df
          13536 => x"7d", -- $034e0
          13537 => x"7f", -- $034e1
          13538 => x"80", -- $034e2
          13539 => x"7f", -- $034e3
          13540 => x"7f", -- $034e4
          13541 => x"7f", -- $034e5
          13542 => x"80", -- $034e6
          13543 => x"81", -- $034e7
          13544 => x"84", -- $034e8
          13545 => x"85", -- $034e9
          13546 => x"84", -- $034ea
          13547 => x"82", -- $034eb
          13548 => x"80", -- $034ec
          13549 => x"80", -- $034ed
          13550 => x"80", -- $034ee
          13551 => x"80", -- $034ef
          13552 => x"7e", -- $034f0
          13553 => x"7c", -- $034f1
          13554 => x"7b", -- $034f2
          13555 => x"7a", -- $034f3
          13556 => x"7a", -- $034f4
          13557 => x"7e", -- $034f5
          13558 => x"80", -- $034f6
          13559 => x"82", -- $034f7
          13560 => x"83", -- $034f8
          13561 => x"84", -- $034f9
          13562 => x"85", -- $034fa
          13563 => x"85", -- $034fb
          13564 => x"86", -- $034fc
          13565 => x"86", -- $034fd
          13566 => x"84", -- $034fe
          13567 => x"81", -- $034ff
          13568 => x"80", -- $03500
          13569 => x"7e", -- $03501
          13570 => x"7c", -- $03502
          13571 => x"7a", -- $03503
          13572 => x"7a", -- $03504
          13573 => x"78", -- $03505
          13574 => x"79", -- $03506
          13575 => x"7b", -- $03507
          13576 => x"7e", -- $03508
          13577 => x"80", -- $03509
          13578 => x"83", -- $0350a
          13579 => x"85", -- $0350b
          13580 => x"85", -- $0350c
          13581 => x"85", -- $0350d
          13582 => x"87", -- $0350e
          13583 => x"88", -- $0350f
          13584 => x"85", -- $03510
          13585 => x"82", -- $03511
          13586 => x"81", -- $03512
          13587 => x"7f", -- $03513
          13588 => x"7f", -- $03514
          13589 => x"80", -- $03515
          13590 => x"80", -- $03516
          13591 => x"80", -- $03517
          13592 => x"7f", -- $03518
          13593 => x"7f", -- $03519
          13594 => x"80", -- $0351a
          13595 => x"80", -- $0351b
          13596 => x"82", -- $0351c
          13597 => x"83", -- $0351d
          13598 => x"82", -- $0351e
          13599 => x"80", -- $0351f
          13600 => x"80", -- $03520
          13601 => x"80", -- $03521
          13602 => x"7f", -- $03522
          13603 => x"7f", -- $03523
          13604 => x"7f", -- $03524
          13605 => x"7d", -- $03525
          13606 => x"7c", -- $03526
          13607 => x"7c", -- $03527
          13608 => x"7d", -- $03528
          13609 => x"7e", -- $03529
          13610 => x"80", -- $0352a
          13611 => x"81", -- $0352b
          13612 => x"82", -- $0352c
          13613 => x"82", -- $0352d
          13614 => x"82", -- $0352e
          13615 => x"83", -- $0352f
          13616 => x"82", -- $03530
          13617 => x"83", -- $03531
          13618 => x"83", -- $03532
          13619 => x"80", -- $03533
          13620 => x"80", -- $03534
          13621 => x"81", -- $03535
          13622 => x"82", -- $03536
          13623 => x"82", -- $03537
          13624 => x"84", -- $03538
          13625 => x"86", -- $03539
          13626 => x"86", -- $0353a
          13627 => x"86", -- $0353b
          13628 => x"86", -- $0353c
          13629 => x"85", -- $0353d
          13630 => x"85", -- $0353e
          13631 => x"84", -- $0353f
          13632 => x"85", -- $03540
          13633 => x"83", -- $03541
          13634 => x"82", -- $03542
          13635 => x"81", -- $03543
          13636 => x"7f", -- $03544
          13637 => x"7d", -- $03545
          13638 => x"7c", -- $03546
          13639 => x"7b", -- $03547
          13640 => x"7a", -- $03548
          13641 => x"79", -- $03549
          13642 => x"79", -- $0354a
          13643 => x"7a", -- $0354b
          13644 => x"7c", -- $0354c
          13645 => x"7e", -- $0354d
          13646 => x"80", -- $0354e
          13647 => x"81", -- $0354f
          13648 => x"84", -- $03550
          13649 => x"86", -- $03551
          13650 => x"87", -- $03552
          13651 => x"88", -- $03553
          13652 => x"88", -- $03554
          13653 => x"88", -- $03555
          13654 => x"87", -- $03556
          13655 => x"85", -- $03557
          13656 => x"82", -- $03558
          13657 => x"80", -- $03559
          13658 => x"7e", -- $0355a
          13659 => x"7b", -- $0355b
          13660 => x"7b", -- $0355c
          13661 => x"7a", -- $0355d
          13662 => x"7a", -- $0355e
          13663 => x"7a", -- $0355f
          13664 => x"7c", -- $03560
          13665 => x"7e", -- $03561
          13666 => x"80", -- $03562
          13667 => x"83", -- $03563
          13668 => x"87", -- $03564
          13669 => x"89", -- $03565
          13670 => x"8a", -- $03566
          13671 => x"8a", -- $03567
          13672 => x"8a", -- $03568
          13673 => x"8a", -- $03569
          13674 => x"88", -- $0356a
          13675 => x"86", -- $0356b
          13676 => x"83", -- $0356c
          13677 => x"80", -- $0356d
          13678 => x"80", -- $0356e
          13679 => x"7e", -- $0356f
          13680 => x"7d", -- $03570
          13681 => x"7c", -- $03571
          13682 => x"7b", -- $03572
          13683 => x"7c", -- $03573
          13684 => x"7e", -- $03574
          13685 => x"7f", -- $03575
          13686 => x"81", -- $03576
          13687 => x"83", -- $03577
          13688 => x"83", -- $03578
          13689 => x"83", -- $03579
          13690 => x"83", -- $0357a
          13691 => x"83", -- $0357b
          13692 => x"82", -- $0357c
          13693 => x"82", -- $0357d
          13694 => x"82", -- $0357e
          13695 => x"81", -- $0357f
          13696 => x"80", -- $03580
          13697 => x"80", -- $03581
          13698 => x"80", -- $03582
          13699 => x"80", -- $03583
          13700 => x"81", -- $03584
          13701 => x"81", -- $03585
          13702 => x"81", -- $03586
          13703 => x"82", -- $03587
          13704 => x"83", -- $03588
          13705 => x"84", -- $03589
          13706 => x"85", -- $0358a
          13707 => x"84", -- $0358b
          13708 => x"83", -- $0358c
          13709 => x"82", -- $0358d
          13710 => x"80", -- $0358e
          13711 => x"80", -- $0358f
          13712 => x"7e", -- $03590
          13713 => x"7c", -- $03591
          13714 => x"7b", -- $03592
          13715 => x"7a", -- $03593
          13716 => x"7a", -- $03594
          13717 => x"7c", -- $03595
          13718 => x"7f", -- $03596
          13719 => x"80", -- $03597
          13720 => x"82", -- $03598
          13721 => x"84", -- $03599
          13722 => x"85", -- $0359a
          13723 => x"86", -- $0359b
          13724 => x"87", -- $0359c
          13725 => x"89", -- $0359d
          13726 => x"89", -- $0359e
          13727 => x"88", -- $0359f
          13728 => x"86", -- $035a0
          13729 => x"86", -- $035a1
          13730 => x"86", -- $035a2
          13731 => x"85", -- $035a3
          13732 => x"86", -- $035a4
          13733 => x"83", -- $035a5
          13734 => x"80", -- $035a6
          13735 => x"80", -- $035a7
          13736 => x"82", -- $035a8
          13737 => x"83", -- $035a9
          13738 => x"83", -- $035aa
          13739 => x"83", -- $035ab
          13740 => x"82", -- $035ac
          13741 => x"81", -- $035ad
          13742 => x"80", -- $035ae
          13743 => x"81", -- $035af
          13744 => x"80", -- $035b0
          13745 => x"7b", -- $035b1
          13746 => x"78", -- $035b2
          13747 => x"77", -- $035b3
          13748 => x"75", -- $035b4
          13749 => x"75", -- $035b5
          13750 => x"77", -- $035b6
          13751 => x"78", -- $035b7
          13752 => x"7a", -- $035b8
          13753 => x"7d", -- $035b9
          13754 => x"81", -- $035ba
          13755 => x"85", -- $035bb
          13756 => x"87", -- $035bc
          13757 => x"8a", -- $035bd
          13758 => x"8b", -- $035be
          13759 => x"89", -- $035bf
          13760 => x"89", -- $035c0
          13761 => x"88", -- $035c1
          13762 => x"85", -- $035c2
          13763 => x"81", -- $035c3
          13764 => x"7d", -- $035c4
          13765 => x"79", -- $035c5
          13766 => x"76", -- $035c6
          13767 => x"75", -- $035c7
          13768 => x"75", -- $035c8
          13769 => x"76", -- $035c9
          13770 => x"78", -- $035ca
          13771 => x"7a", -- $035cb
          13772 => x"7f", -- $035cc
          13773 => x"82", -- $035cd
          13774 => x"87", -- $035ce
          13775 => x"8a", -- $035cf
          13776 => x"8c", -- $035d0
          13777 => x"8e", -- $035d1
          13778 => x"8d", -- $035d2
          13779 => x"8c", -- $035d3
          13780 => x"89", -- $035d4
          13781 => x"86", -- $035d5
          13782 => x"84", -- $035d6
          13783 => x"80", -- $035d7
          13784 => x"7f", -- $035d8
          13785 => x"7c", -- $035d9
          13786 => x"7c", -- $035da
          13787 => x"7b", -- $035db
          13788 => x"7e", -- $035dc
          13789 => x"80", -- $035dd
          13790 => x"81", -- $035de
          13791 => x"83", -- $035df
          13792 => x"86", -- $035e0
          13793 => x"87", -- $035e1
          13794 => x"87", -- $035e2
          13795 => x"88", -- $035e3
          13796 => x"87", -- $035e4
          13797 => x"84", -- $035e5
          13798 => x"80", -- $035e6
          13799 => x"7e", -- $035e7
          13800 => x"7c", -- $035e8
          13801 => x"79", -- $035e9
          13802 => x"77", -- $035ea
          13803 => x"76", -- $035eb
          13804 => x"75", -- $035ec
          13805 => x"77", -- $035ed
          13806 => x"79", -- $035ee
          13807 => x"7c", -- $035ef
          13808 => x"7e", -- $035f0
          13809 => x"80", -- $035f1
          13810 => x"81", -- $035f2
          13811 => x"82", -- $035f3
          13812 => x"83", -- $035f4
          13813 => x"83", -- $035f5
          13814 => x"83", -- $035f6
          13815 => x"80", -- $035f7
          13816 => x"7f", -- $035f8
          13817 => x"7f", -- $035f9
          13818 => x"7e", -- $035fa
          13819 => x"7e", -- $035fb
          13820 => x"7e", -- $035fc
          13821 => x"7f", -- $035fd
          13822 => x"7f", -- $035fe
          13823 => x"80", -- $035ff
          13824 => x"84", -- $03600
          13825 => x"86", -- $03601
          13826 => x"88", -- $03602
          13827 => x"8a", -- $03603
          13828 => x"8a", -- $03604
          13829 => x"8b", -- $03605
          13830 => x"8b", -- $03606
          13831 => x"8c", -- $03607
          13832 => x"8a", -- $03608
          13833 => x"88", -- $03609
          13834 => x"86", -- $0360a
          13835 => x"85", -- $0360b
          13836 => x"85", -- $0360c
          13837 => x"82", -- $0360d
          13838 => x"7e", -- $0360e
          13839 => x"7e", -- $0360f
          13840 => x"7f", -- $03610
          13841 => x"80", -- $03611
          13842 => x"81", -- $03612
          13843 => x"81", -- $03613
          13844 => x"81", -- $03614
          13845 => x"7f", -- $03615
          13846 => x"80", -- $03616
          13847 => x"81", -- $03617
          13848 => x"7f", -- $03618
          13849 => x"7c", -- $03619
          13850 => x"79", -- $0361a
          13851 => x"77", -- $0361b
          13852 => x"76", -- $0361c
          13853 => x"77", -- $0361d
          13854 => x"78", -- $0361e
          13855 => x"79", -- $0361f
          13856 => x"79", -- $03620
          13857 => x"7d", -- $03621
          13858 => x"80", -- $03622
          13859 => x"83", -- $03623
          13860 => x"87", -- $03624
          13861 => x"88", -- $03625
          13862 => x"88", -- $03626
          13863 => x"88", -- $03627
          13864 => x"8a", -- $03628
          13865 => x"88", -- $03629
          13866 => x"84", -- $0362a
          13867 => x"80", -- $0362b
          13868 => x"7d", -- $0362c
          13869 => x"79", -- $0362d
          13870 => x"78", -- $0362e
          13871 => x"77", -- $0362f
          13872 => x"76", -- $03630
          13873 => x"76", -- $03631
          13874 => x"78", -- $03632
          13875 => x"7b", -- $03633
          13876 => x"7f", -- $03634
          13877 => x"82", -- $03635
          13878 => x"86", -- $03636
          13879 => x"88", -- $03637
          13880 => x"8a", -- $03638
          13881 => x"8c", -- $03639
          13882 => x"8d", -- $0363a
          13883 => x"8d", -- $0363b
          13884 => x"8b", -- $0363c
          13885 => x"88", -- $0363d
          13886 => x"83", -- $0363e
          13887 => x"80", -- $0363f
          13888 => x"80", -- $03640
          13889 => x"7e", -- $03641
          13890 => x"7d", -- $03642
          13891 => x"7c", -- $03643
          13892 => x"7c", -- $03644
          13893 => x"7d", -- $03645
          13894 => x"80", -- $03646
          13895 => x"83", -- $03647
          13896 => x"84", -- $03648
          13897 => x"85", -- $03649
          13898 => x"85", -- $0364a
          13899 => x"85", -- $0364b
          13900 => x"85", -- $0364c
          13901 => x"84", -- $0364d
          13902 => x"82", -- $0364e
          13903 => x"7f", -- $0364f
          13904 => x"7b", -- $03650
          13905 => x"7a", -- $03651
          13906 => x"79", -- $03652
          13907 => x"79", -- $03653
          13908 => x"79", -- $03654
          13909 => x"79", -- $03655
          13910 => x"79", -- $03656
          13911 => x"7b", -- $03657
          13912 => x"7e", -- $03658
          13913 => x"80", -- $03659
          13914 => x"80", -- $0365a
          13915 => x"80", -- $0365b
          13916 => x"80", -- $0365c
          13917 => x"80", -- $0365d
          13918 => x"80", -- $0365e
          13919 => x"80", -- $0365f
          13920 => x"7f", -- $03660
          13921 => x"7d", -- $03661
          13922 => x"7d", -- $03662
          13923 => x"7d", -- $03663
          13924 => x"7d", -- $03664
          13925 => x"7d", -- $03665
          13926 => x"7d", -- $03666
          13927 => x"7f", -- $03667
          13928 => x"81", -- $03668
          13929 => x"84", -- $03669
          13930 => x"87", -- $0366a
          13931 => x"88", -- $0366b
          13932 => x"88", -- $0366c
          13933 => x"8a", -- $0366d
          13934 => x"8b", -- $0366e
          13935 => x"8a", -- $0366f
          13936 => x"89", -- $03670
          13937 => x"86", -- $03671
          13938 => x"84", -- $03672
          13939 => x"83", -- $03673
          13940 => x"82", -- $03674
          13941 => x"81", -- $03675
          13942 => x"80", -- $03676
          13943 => x"80", -- $03677
          13944 => x"80", -- $03678
          13945 => x"80", -- $03679
          13946 => x"80", -- $0367a
          13947 => x"80", -- $0367b
          13948 => x"80", -- $0367c
          13949 => x"7f", -- $0367d
          13950 => x"7f", -- $0367e
          13951 => x"7f", -- $0367f
          13952 => x"7e", -- $03680
          13953 => x"7c", -- $03681
          13954 => x"7a", -- $03682
          13955 => x"78", -- $03683
          13956 => x"77", -- $03684
          13957 => x"77", -- $03685
          13958 => x"78", -- $03686
          13959 => x"78", -- $03687
          13960 => x"78", -- $03688
          13961 => x"7a", -- $03689
          13962 => x"7c", -- $0368a
          13963 => x"7e", -- $0368b
          13964 => x"7f", -- $0368c
          13965 => x"80", -- $0368d
          13966 => x"80", -- $0368e
          13967 => x"81", -- $0368f
          13968 => x"82", -- $03690
          13969 => x"83", -- $03691
          13970 => x"82", -- $03692
          13971 => x"81", -- $03693
          13972 => x"80", -- $03694
          13973 => x"7f", -- $03695
          13974 => x"7f", -- $03696
          13975 => x"7f", -- $03697
          13976 => x"7f", -- $03698
          13977 => x"7e", -- $03699
          13978 => x"80", -- $0369a
          13979 => x"80", -- $0369b
          13980 => x"82", -- $0369c
          13981 => x"84", -- $0369d
          13982 => x"85", -- $0369e
          13983 => x"85", -- $0369f
          13984 => x"86", -- $036a0
          13985 => x"88", -- $036a1
          13986 => x"88", -- $036a2
          13987 => x"87", -- $036a3
          13988 => x"86", -- $036a4
          13989 => x"84", -- $036a5
          13990 => x"83", -- $036a6
          13991 => x"82", -- $036a7
          13992 => x"81", -- $036a8
          13993 => x"80", -- $036a9
          13994 => x"7d", -- $036aa
          13995 => x"7c", -- $036ab
          13996 => x"7c", -- $036ac
          13997 => x"7c", -- $036ad
          13998 => x"7b", -- $036ae
          13999 => x"7a", -- $036af
          14000 => x"7a", -- $036b0
          14001 => x"7a", -- $036b1
          14002 => x"7b", -- $036b2
          14003 => x"7b", -- $036b3
          14004 => x"7a", -- $036b4
          14005 => x"79", -- $036b5
          14006 => x"79", -- $036b6
          14007 => x"7a", -- $036b7
          14008 => x"7a", -- $036b8
          14009 => x"7b", -- $036b9
          14010 => x"7b", -- $036ba
          14011 => x"7b", -- $036bb
          14012 => x"7c", -- $036bc
          14013 => x"7d", -- $036bd
          14014 => x"7e", -- $036be
          14015 => x"7e", -- $036bf
          14016 => x"7f", -- $036c0
          14017 => x"80", -- $036c1
          14018 => x"80", -- $036c2
          14019 => x"81", -- $036c3
          14020 => x"81", -- $036c4
          14021 => x"80", -- $036c5
          14022 => x"80", -- $036c6
          14023 => x"80", -- $036c7
          14024 => x"80", -- $036c8
          14025 => x"80", -- $036c9
          14026 => x"7f", -- $036ca
          14027 => x"7f", -- $036cb
          14028 => x"7f", -- $036cc
          14029 => x"7f", -- $036cd
          14030 => x"80", -- $036ce
          14031 => x"7f", -- $036cf
          14032 => x"80", -- $036d0
          14033 => x"80", -- $036d1
          14034 => x"80", -- $036d2
          14035 => x"81", -- $036d3
          14036 => x"82", -- $036d4
          14037 => x"82", -- $036d5
          14038 => x"82", -- $036d6
          14039 => x"82", -- $036d7
          14040 => x"83", -- $036d8
          14041 => x"83", -- $036d9
          14042 => x"82", -- $036da
          14043 => x"81", -- $036db
          14044 => x"80", -- $036dc
          14045 => x"80", -- $036dd
          14046 => x"80", -- $036de
          14047 => x"7f", -- $036df
          14048 => x"7e", -- $036e0
          14049 => x"7d", -- $036e1
          14050 => x"7d", -- $036e2
          14051 => x"7d", -- $036e3
          14052 => x"7d", -- $036e4
          14053 => x"7c", -- $036e5
          14054 => x"7c", -- $036e6
          14055 => x"7c", -- $036e7
          14056 => x"7c", -- $036e8
          14057 => x"7d", -- $036e9
          14058 => x"7d", -- $036ea
          14059 => x"7d", -- $036eb
          14060 => x"7d", -- $036ec
          14061 => x"7e", -- $036ed
          14062 => x"7e", -- $036ee
          14063 => x"7f", -- $036ef
          14064 => x"7f", -- $036f0
          14065 => x"7f", -- $036f1
          14066 => x"80", -- $036f2
          14067 => x"80", -- $036f3
          14068 => x"80", -- $036f4
          14069 => x"80", -- $036f5
          14070 => x"80", -- $036f6
          14071 => x"80", -- $036f7
          14072 => x"80", -- $036f8
          14073 => x"80", -- $036f9
          14074 => x"80", -- $036fa
          14075 => x"80", -- $036fb
          14076 => x"80", -- $036fc
          14077 => x"7f", -- $036fd
          14078 => x"7e", -- $036fe
          14079 => x"7e", -- $036ff
          14080 => x"7d", -- $03700
          14081 => x"7d", -- $03701
          14082 => x"7d", -- $03702
          14083 => x"7d", -- $03703
          14084 => x"7d", -- $03704
          14085 => x"7e", -- $03705
          14086 => x"7f", -- $03706
          14087 => x"80", -- $03707
          14088 => x"80", -- $03708
          14089 => x"80", -- $03709
          14090 => x"80", -- $0370a
          14091 => x"81", -- $0370b
          14092 => x"81", -- $0370c
          14093 => x"81", -- $0370d
          14094 => x"81", -- $0370e
          14095 => x"81", -- $0370f
          14096 => x"81", -- $03710
          14097 => x"80", -- $03711
          14098 => x"80", -- $03712
          14099 => x"80", -- $03713
          14100 => x"80", -- $03714
          14101 => x"80", -- $03715
          14102 => x"80", -- $03716
          14103 => x"7f", -- $03717
          14104 => x"7f", -- $03718
          14105 => x"7e", -- $03719
          14106 => x"7f", -- $0371a
          14107 => x"7e", -- $0371b
          14108 => x"7e", -- $0371c
          14109 => x"7e", -- $0371d
          14110 => x"7e", -- $0371e
          14111 => x"7e", -- $0371f
          14112 => x"7f", -- $03720
          14113 => x"7f", -- $03721
          14114 => x"7f", -- $03722
          14115 => x"7f", -- $03723
          14116 => x"7f", -- $03724
          14117 => x"80", -- $03725
          14118 => x"80", -- $03726
          14119 => x"80", -- $03727
          14120 => x"80", -- $03728
          14121 => x"80", -- $03729
          14122 => x"80", -- $0372a
          14123 => x"80", -- $0372b
          14124 => x"80", -- $0372c
          14125 => x"80", -- $0372d
          14126 => x"80", -- $0372e
          14127 => x"80", -- $0372f
          14128 => x"80", -- $03730
          14129 => x"80", -- $03731
          14130 => x"7f", -- $03732
          14131 => x"7f", -- $03733
          14132 => x"7f", -- $03734
          14133 => x"7f", -- $03735
          14134 => x"7f", -- $03736
          14135 => x"7f", -- $03737
          14136 => x"7f", -- $03738
          14137 => x"7f", -- $03739
          14138 => x"80", -- $0373a
          14139 => x"80", -- $0373b
          14140 => x"80", -- $0373c
          14141 => x"80", -- $0373d
          14142 => x"80", -- $0373e
          14143 => x"80", -- $0373f
          14144 => x"80", -- $03740
          14145 => x"80", -- $03741
          14146 => x"80", -- $03742
          14147 => x"80", -- $03743
          14148 => x"7e", -- $03744
          14149 => x"7e", -- $03745
          14150 => x"7e", -- $03746
          14151 => x"7e", -- $03747
          14152 => x"7c", -- $03748
          14153 => x"7b", -- $03749
          14154 => x"7b", -- $0374a
          14155 => x"7c", -- $0374b
          14156 => x"7c", -- $0374c
          14157 => x"7b", -- $0374d
          14158 => x"7b", -- $0374e
          14159 => x"7b", -- $0374f
          14160 => x"7c", -- $03750
          14161 => x"7d", -- $03751
          14162 => x"7d", -- $03752
          14163 => x"7d", -- $03753
          14164 => x"7e", -- $03754
          14165 => x"7f", -- $03755
          14166 => x"7f", -- $03756
          14167 => x"80", -- $03757
          14168 => x"7f", -- $03758
          14169 => x"7f", -- $03759
          14170 => x"80", -- $0375a
          14171 => x"80", -- $0375b
          14172 => x"81", -- $0375c
          14173 => x"81", -- $0375d
          14174 => x"81", -- $0375e
          14175 => x"82", -- $0375f
          14176 => x"83", -- $03760
          14177 => x"83", -- $03761
          14178 => x"83", -- $03762
          14179 => x"83", -- $03763
          14180 => x"82", -- $03764
          14181 => x"82", -- $03765
          14182 => x"80", -- $03766
          14183 => x"80", -- $03767
          14184 => x"80", -- $03768
          14185 => x"7f", -- $03769
          14186 => x"7e", -- $0376a
          14187 => x"7e", -- $0376b
          14188 => x"7e", -- $0376c
          14189 => x"7e", -- $0376d
          14190 => x"7e", -- $0376e
          14191 => x"7d", -- $0376f
          14192 => x"7d", -- $03770
          14193 => x"7e", -- $03771
          14194 => x"7f", -- $03772
          14195 => x"7f", -- $03773
          14196 => x"7f", -- $03774
          14197 => x"7e", -- $03775
          14198 => x"7f", -- $03776
          14199 => x"7f", -- $03777
          14200 => x"7f", -- $03778
          14201 => x"7d", -- $03779
          14202 => x"7d", -- $0377a
          14203 => x"7d", -- $0377b
          14204 => x"7e", -- $0377c
          14205 => x"7d", -- $0377d
          14206 => x"7b", -- $0377e
          14207 => x"7b", -- $0377f
          14208 => x"7c", -- $03780
          14209 => x"7c", -- $03781
          14210 => x"7b", -- $03782
          14211 => x"7b", -- $03783
          14212 => x"7d", -- $03784
          14213 => x"7e", -- $03785
          14214 => x"7e", -- $03786
          14215 => x"7e", -- $03787
          14216 => x"7f", -- $03788
          14217 => x"80", -- $03789
          14218 => x"80", -- $0378a
          14219 => x"7f", -- $0378b
          14220 => x"80", -- $0378c
          14221 => x"80", -- $0378d
          14222 => x"80", -- $0378e
          14223 => x"80", -- $0378f
          14224 => x"80", -- $03790
          14225 => x"80", -- $03791
          14226 => x"80", -- $03792
          14227 => x"80", -- $03793
          14228 => x"80", -- $03794
          14229 => x"80", -- $03795
          14230 => x"80", -- $03796
          14231 => x"80", -- $03797
          14232 => x"80", -- $03798
          14233 => x"80", -- $03799
          14234 => x"80", -- $0379a
          14235 => x"7f", -- $0379b
          14236 => x"80", -- $0379c
          14237 => x"7f", -- $0379d
          14238 => x"7e", -- $0379e
          14239 => x"7e", -- $0379f
          14240 => x"7e", -- $037a0
          14241 => x"7f", -- $037a1
          14242 => x"7f", -- $037a2
          14243 => x"7f", -- $037a3
          14244 => x"7f", -- $037a4
          14245 => x"80", -- $037a5
          14246 => x"80", -- $037a6
          14247 => x"80", -- $037a7
          14248 => x"80", -- $037a8
          14249 => x"80", -- $037a9
          14250 => x"81", -- $037aa
          14251 => x"80", -- $037ab
          14252 => x"80", -- $037ac
          14253 => x"80", -- $037ad
          14254 => x"80", -- $037ae
          14255 => x"80", -- $037af
          14256 => x"7f", -- $037b0
          14257 => x"7f", -- $037b1
          14258 => x"7f", -- $037b2
          14259 => x"7e", -- $037b3
          14260 => x"7e", -- $037b4
          14261 => x"7d", -- $037b5
          14262 => x"7e", -- $037b6
          14263 => x"7e", -- $037b7
          14264 => x"7e", -- $037b8
          14265 => x"7f", -- $037b9
          14266 => x"7f", -- $037ba
          14267 => x"7f", -- $037bb
          14268 => x"7f", -- $037bc
          14269 => x"7f", -- $037bd
          14270 => x"7f", -- $037be
          14271 => x"80", -- $037bf
          14272 => x"80", -- $037c0
          14273 => x"7f", -- $037c1
          14274 => x"7f", -- $037c2
          14275 => x"7f", -- $037c3
          14276 => x"80", -- $037c4
          14277 => x"80", -- $037c5
          14278 => x"80", -- $037c6
          14279 => x"80", -- $037c7
          14280 => x"80", -- $037c8
          14281 => x"80", -- $037c9
          14282 => x"80", -- $037ca
          14283 => x"80", -- $037cb
          14284 => x"80", -- $037cc
          14285 => x"80", -- $037cd
          14286 => x"81", -- $037ce
          14287 => x"81", -- $037cf
          14288 => x"80", -- $037d0
          14289 => x"80", -- $037d1
          14290 => x"80", -- $037d2
          14291 => x"80", -- $037d3
          14292 => x"80", -- $037d4
          14293 => x"80", -- $037d5
          14294 => x"80", -- $037d6
          14295 => x"80", -- $037d7
          14296 => x"80", -- $037d8
          14297 => x"81", -- $037d9
          14298 => x"81", -- $037da
          14299 => x"81", -- $037db
          14300 => x"81", -- $037dc
          14301 => x"81", -- $037dd
          14302 => x"81", -- $037de
          14303 => x"81", -- $037df
          14304 => x"81", -- $037e0
          14305 => x"81", -- $037e1
          14306 => x"81", -- $037e2
          14307 => x"81", -- $037e3
          14308 => x"80", -- $037e4
          14309 => x"80", -- $037e5
          14310 => x"80", -- $037e6
          14311 => x"80", -- $037e7
          14312 => x"7f", -- $037e8
          14313 => x"7f", -- $037e9
          14314 => x"80", -- $037ea
          14315 => x"80", -- $037eb
          14316 => x"7f", -- $037ec
          14317 => x"80", -- $037ed
          14318 => x"80", -- $037ee
          14319 => x"80", -- $037ef
          14320 => x"80", -- $037f0
          14321 => x"80", -- $037f1
          14322 => x"80", -- $037f2
          14323 => x"80", -- $037f3
          14324 => x"80", -- $037f4
          14325 => x"80", -- $037f5
          14326 => x"80", -- $037f6
          14327 => x"80", -- $037f7
          14328 => x"80", -- $037f8
          14329 => x"80", -- $037f9
          14330 => x"80", -- $037fa
          14331 => x"81", -- $037fb
          14332 => x"80", -- $037fc
          14333 => x"81", -- $037fd
          14334 => x"80", -- $037fe
          14335 => x"81", -- $037ff
          14336 => x"80", -- $03800
          14337 => x"80", -- $03801
          14338 => x"80", -- $03802
          14339 => x"80", -- $03803
          14340 => x"80", -- $03804
          14341 => x"7f", -- $03805
          14342 => x"80", -- $03806
          14343 => x"80", -- $03807
          14344 => x"80", -- $03808
          14345 => x"80", -- $03809
          14346 => x"80", -- $0380a
          14347 => x"80", -- $0380b
          14348 => x"80", -- $0380c
          14349 => x"80", -- $0380d
          14350 => x"80", -- $0380e
          14351 => x"81", -- $0380f
          14352 => x"80", -- $03810
          14353 => x"80", -- $03811
          14354 => x"81", -- $03812
          14355 => x"81", -- $03813
          14356 => x"80", -- $03814
          14357 => x"80", -- $03815
          14358 => x"81", -- $03816
          14359 => x"80", -- $03817
          14360 => x"80", -- $03818
          14361 => x"80", -- $03819
          14362 => x"80", -- $0381a
          14363 => x"81", -- $0381b
          14364 => x"80", -- $0381c
          14365 => x"80", -- $0381d
          14366 => x"80", -- $0381e
          14367 => x"80", -- $0381f
          14368 => x"81", -- $03820
          14369 => x"81", -- $03821
          14370 => x"81", -- $03822
          14371 => x"81", -- $03823
          14372 => x"82", -- $03824
          14373 => x"82", -- $03825
          14374 => x"80", -- $03826
          14375 => x"80", -- $03827
          14376 => x"81", -- $03828
          14377 => x"80", -- $03829
          14378 => x"80", -- $0382a
          14379 => x"80", -- $0382b
          14380 => x"81", -- $0382c
          14381 => x"80", -- $0382d
          14382 => x"80", -- $0382e
          14383 => x"80", -- $0382f
          14384 => x"81", -- $03830
          14385 => x"80", -- $03831
          14386 => x"80", -- $03832
          14387 => x"80", -- $03833
          14388 => x"80", -- $03834
          14389 => x"80", -- $03835
          14390 => x"7f", -- $03836
          14391 => x"7f", -- $03837
          14392 => x"7f", -- $03838
          14393 => x"7f", -- $03839
          14394 => x"7f", -- $0383a
          14395 => x"7f", -- $0383b
          14396 => x"7f", -- $0383c
          14397 => x"7f", -- $0383d
          14398 => x"7f", -- $0383e
          14399 => x"80", -- $0383f
          14400 => x"80", -- $03840
          14401 => x"80", -- $03841
          14402 => x"80", -- $03842
          14403 => x"81", -- $03843
          14404 => x"81", -- $03844
          14405 => x"81", -- $03845
          14406 => x"81", -- $03846
          14407 => x"81", -- $03847
          14408 => x"81", -- $03848
          14409 => x"81", -- $03849
          14410 => x"81", -- $0384a
          14411 => x"81", -- $0384b
          14412 => x"81", -- $0384c
          14413 => x"81", -- $0384d
          14414 => x"80", -- $0384e
          14415 => x"81", -- $0384f
          14416 => x"81", -- $03850
          14417 => x"81", -- $03851
          14418 => x"81", -- $03852
          14419 => x"82", -- $03853
          14420 => x"81", -- $03854
          14421 => x"81", -- $03855
          14422 => x"81", -- $03856
          14423 => x"81", -- $03857
          14424 => x"81", -- $03858
          14425 => x"81", -- $03859
          14426 => x"80", -- $0385a
          14427 => x"80", -- $0385b
          14428 => x"80", -- $0385c
          14429 => x"80", -- $0385d
          14430 => x"80", -- $0385e
          14431 => x"80", -- $0385f
          14432 => x"80", -- $03860
          14433 => x"80", -- $03861
          14434 => x"80", -- $03862
          14435 => x"80", -- $03863
          14436 => x"80", -- $03864
          14437 => x"80", -- $03865
          14438 => x"81", -- $03866
          14439 => x"81", -- $03867
          14440 => x"80", -- $03868
          14441 => x"80", -- $03869
          14442 => x"80", -- $0386a
          14443 => x"80", -- $0386b
          14444 => x"80", -- $0386c
          14445 => x"80", -- $0386d
          14446 => x"80", -- $0386e
          14447 => x"80", -- $0386f
          14448 => x"80", -- $03870
          14449 => x"80", -- $03871
          14450 => x"81", -- $03872
          14451 => x"81", -- $03873
          14452 => x"80", -- $03874
          14453 => x"81", -- $03875
          14454 => x"81", -- $03876
          14455 => x"81", -- $03877
          14456 => x"81", -- $03878
          14457 => x"81", -- $03879
          14458 => x"81", -- $0387a
          14459 => x"81", -- $0387b
          14460 => x"80", -- $0387c
          14461 => x"81", -- $0387d
          14462 => x"81", -- $0387e
          14463 => x"80", -- $0387f
          14464 => x"80", -- $03880
          14465 => x"80", -- $03881
          14466 => x"80", -- $03882
          14467 => x"80", -- $03883
          14468 => x"80", -- $03884
          14469 => x"80", -- $03885
          14470 => x"81", -- $03886
          14471 => x"81", -- $03887
          14472 => x"81", -- $03888
          14473 => x"81", -- $03889
          14474 => x"80", -- $0388a
          14475 => x"81", -- $0388b
          14476 => x"81", -- $0388c
          14477 => x"81", -- $0388d
          14478 => x"81", -- $0388e
          14479 => x"81", -- $0388f
          14480 => x"81", -- $03890
          14481 => x"81", -- $03891
          14482 => x"81", -- $03892
          14483 => x"82", -- $03893
          14484 => x"80", -- $03894
          14485 => x"81", -- $03895
          14486 => x"83", -- $03896
          14487 => x"82", -- $03897
          14488 => x"81", -- $03898
          14489 => x"83", -- $03899
          14490 => x"82", -- $0389a
          14491 => x"82", -- $0389b
          14492 => x"82", -- $0389c
          14493 => x"82", -- $0389d
          14494 => x"81", -- $0389e
          14495 => x"81", -- $0389f
          14496 => x"81", -- $038a0
          14497 => x"81", -- $038a1
          14498 => x"81", -- $038a2
          14499 => x"80", -- $038a3
          14500 => x"81", -- $038a4
          14501 => x"81", -- $038a5
          14502 => x"80", -- $038a6
          14503 => x"81", -- $038a7
          14504 => x"81", -- $038a8
          14505 => x"80", -- $038a9
          14506 => x"80", -- $038aa
          14507 => x"81", -- $038ab
          14508 => x"81", -- $038ac
          14509 => x"81", -- $038ad
          14510 => x"81", -- $038ae
          14511 => x"80", -- $038af
          14512 => x"81", -- $038b0
          14513 => x"80", -- $038b1
          14514 => x"80", -- $038b2
          14515 => x"81", -- $038b3
          14516 => x"80", -- $038b4
          14517 => x"80", -- $038b5
          14518 => x"80", -- $038b6
          14519 => x"80", -- $038b7
          14520 => x"82", -- $038b8
          14521 => x"81", -- $038b9
          14522 => x"81", -- $038ba
          14523 => x"82", -- $038bb
          14524 => x"81", -- $038bc
          14525 => x"81", -- $038bd
          14526 => x"82", -- $038be
          14527 => x"82", -- $038bf
          14528 => x"81", -- $038c0
          14529 => x"81", -- $038c1
          14530 => x"82", -- $038c2
          14531 => x"81", -- $038c3
          14532 => x"81", -- $038c4
          14533 => x"82", -- $038c5
          14534 => x"82", -- $038c6
          14535 => x"81", -- $038c7
          14536 => x"82", -- $038c8
          14537 => x"81", -- $038c9
          14538 => x"81", -- $038ca
          14539 => x"82", -- $038cb
          14540 => x"81", -- $038cc
          14541 => x"81", -- $038cd
          14542 => x"82", -- $038ce
          14543 => x"81", -- $038cf
          14544 => x"82", -- $038d0
          14545 => x"81", -- $038d1
          14546 => x"81", -- $038d2
          14547 => x"81", -- $038d3
          14548 => x"80", -- $038d4
          14549 => x"81", -- $038d5
          14550 => x"81", -- $038d6
          14551 => x"82", -- $038d7
          14552 => x"80", -- $038d8
          14553 => x"80", -- $038d9
          14554 => x"82", -- $038da
          14555 => x"81", -- $038db
          14556 => x"81", -- $038dc
          14557 => x"81", -- $038dd
          14558 => x"82", -- $038de
          14559 => x"82", -- $038df
          14560 => x"81", -- $038e0
          14561 => x"82", -- $038e1
          14562 => x"81", -- $038e2
          14563 => x"81", -- $038e3
          14564 => x"81", -- $038e4
          14565 => x"81", -- $038e5
          14566 => x"81", -- $038e6
          14567 => x"81", -- $038e7
          14568 => x"81", -- $038e8
          14569 => x"81", -- $038e9
          14570 => x"80", -- $038ea
          14571 => x"80", -- $038eb
          14572 => x"81", -- $038ec
          14573 => x"81", -- $038ed
          14574 => x"81", -- $038ee
          14575 => x"81", -- $038ef
          14576 => x"81", -- $038f0
          14577 => x"81", -- $038f1
          14578 => x"80", -- $038f2
          14579 => x"81", -- $038f3
          14580 => x"80", -- $038f4
          14581 => x"81", -- $038f5
          14582 => x"81", -- $038f6
          14583 => x"80", -- $038f7
          14584 => x"80", -- $038f8
          14585 => x"80", -- $038f9
          14586 => x"81", -- $038fa
          14587 => x"80", -- $038fb
          14588 => x"80", -- $038fc
          14589 => x"81", -- $038fd
          14590 => x"81", -- $038fe
          14591 => x"81", -- $038ff
          14592 => x"81", -- $03900
          14593 => x"82", -- $03901
          14594 => x"81", -- $03902
          14595 => x"81", -- $03903
          14596 => x"82", -- $03904
          14597 => x"81", -- $03905
          14598 => x"81", -- $03906
          14599 => x"81", -- $03907
          14600 => x"81", -- $03908
          14601 => x"81", -- $03909
          14602 => x"80", -- $0390a
          14603 => x"80", -- $0390b
          14604 => x"80", -- $0390c
          14605 => x"81", -- $0390d
          14606 => x"81", -- $0390e
          14607 => x"81", -- $0390f
          14608 => x"81", -- $03910
          14609 => x"81", -- $03911
          14610 => x"81", -- $03912
          14611 => x"81", -- $03913
          14612 => x"81", -- $03914
          14613 => x"81", -- $03915
          14614 => x"81", -- $03916
          14615 => x"81", -- $03917
          14616 => x"81", -- $03918
          14617 => x"81", -- $03919
          14618 => x"80", -- $0391a
          14619 => x"80", -- $0391b
          14620 => x"80", -- $0391c
          14621 => x"80", -- $0391d
          14622 => x"80", -- $0391e
          14623 => x"81", -- $0391f
          14624 => x"80", -- $03920
          14625 => x"80", -- $03921
          14626 => x"80", -- $03922
          14627 => x"80", -- $03923
          14628 => x"80", -- $03924
          14629 => x"80", -- $03925
          14630 => x"80", -- $03926
          14631 => x"80", -- $03927
          14632 => x"80", -- $03928
          14633 => x"80", -- $03929
          14634 => x"80", -- $0392a
          14635 => x"80", -- $0392b
          14636 => x"80", -- $0392c
          14637 => x"80", -- $0392d
          14638 => x"80", -- $0392e
          14639 => x"80", -- $0392f
          14640 => x"80", -- $03930
          14641 => x"80", -- $03931
          14642 => x"80", -- $03932
          14643 => x"80", -- $03933
          14644 => x"81", -- $03934
          14645 => x"81", -- $03935
          14646 => x"81", -- $03936
          14647 => x"80", -- $03937
          14648 => x"81", -- $03938
          14649 => x"80", -- $03939
          14650 => x"80", -- $0393a
          14651 => x"80", -- $0393b
          14652 => x"80", -- $0393c
          14653 => x"80", -- $0393d
          14654 => x"80", -- $0393e
          14655 => x"80", -- $0393f
          14656 => x"80", -- $03940
          14657 => x"80", -- $03941
          14658 => x"80", -- $03942
          14659 => x"80", -- $03943
          14660 => x"80", -- $03944
          14661 => x"80", -- $03945
          14662 => x"80", -- $03946
          14663 => x"80", -- $03947
          14664 => x"80", -- $03948
          14665 => x"80", -- $03949
          14666 => x"80", -- $0394a
          14667 => x"80", -- $0394b
          14668 => x"80", -- $0394c
          14669 => x"80", -- $0394d
          14670 => x"80", -- $0394e
          14671 => x"80", -- $0394f
          14672 => x"80", -- $03950
          14673 => x"80", -- $03951
          14674 => x"80", -- $03952
          14675 => x"80", -- $03953
          14676 => x"80", -- $03954
          14677 => x"80", -- $03955
          14678 => x"80", -- $03956
          14679 => x"80", -- $03957
          14680 => x"81", -- $03958
          14681 => x"81", -- $03959
          14682 => x"80", -- $0395a
          14683 => x"81", -- $0395b
          14684 => x"81", -- $0395c
          14685 => x"80", -- $0395d
          14686 => x"80", -- $0395e
          14687 => x"80", -- $0395f
          14688 => x"80", -- $03960
          14689 => x"80", -- $03961
          14690 => x"80", -- $03962
          14691 => x"80", -- $03963
          14692 => x"80", -- $03964
          14693 => x"80", -- $03965
          14694 => x"80", -- $03966
          14695 => x"80", -- $03967
          14696 => x"80", -- $03968
          14697 => x"80", -- $03969
          14698 => x"80", -- $0396a
          14699 => x"80", -- $0396b
          14700 => x"80", -- $0396c
          14701 => x"80", -- $0396d
          14702 => x"80", -- $0396e
          14703 => x"80", -- $0396f
          14704 => x"7f", -- $03970
          14705 => x"80", -- $03971
          14706 => x"80", -- $03972
          14707 => x"80", -- $03973
          14708 => x"7f", -- $03974
          14709 => x"7f", -- $03975
          14710 => x"7f", -- $03976
          14711 => x"7f", -- $03977
          14712 => x"7f", -- $03978
          14713 => x"7f", -- $03979
          14714 => x"80", -- $0397a
          14715 => x"80", -- $0397b
          14716 => x"80", -- $0397c
          14717 => x"80", -- $0397d
          14718 => x"80", -- $0397e
          14719 => x"80", -- $0397f
          14720 => x"80", -- $03980
          14721 => x"81", -- $03981
          14722 => x"81", -- $03982
          14723 => x"81", -- $03983
          14724 => x"82", -- $03984
          14725 => x"82", -- $03985
          14726 => x"82", -- $03986
          14727 => x"81", -- $03987
          14728 => x"81", -- $03988
          14729 => x"82", -- $03989
          14730 => x"81", -- $0398a
          14731 => x"82", -- $0398b
          14732 => x"82", -- $0398c
          14733 => x"81", -- $0398d
          14734 => x"81", -- $0398e
          14735 => x"81", -- $0398f
          14736 => x"81", -- $03990
          14737 => x"81", -- $03991
          14738 => x"80", -- $03992
          14739 => x"81", -- $03993
          14740 => x"80", -- $03994
          14741 => x"80", -- $03995
          14742 => x"80", -- $03996
          14743 => x"80", -- $03997
          14744 => x"7e", -- $03998
          14745 => x"7e", -- $03999
          14746 => x"7e", -- $0399a
          14747 => x"7e", -- $0399b
          14748 => x"7d", -- $0399c
          14749 => x"7d", -- $0399d
          14750 => x"7d", -- $0399e
          14751 => x"7d", -- $0399f
          14752 => x"7d", -- $039a0
          14753 => x"7d", -- $039a1
          14754 => x"7d", -- $039a2
          14755 => x"7d", -- $039a3
          14756 => x"7d", -- $039a4
          14757 => x"7e", -- $039a5
          14758 => x"7e", -- $039a6
          14759 => x"7f", -- $039a7
          14760 => x"80", -- $039a8
          14761 => x"80", -- $039a9
          14762 => x"80", -- $039aa
          14763 => x"82", -- $039ab
          14764 => x"83", -- $039ac
          14765 => x"83", -- $039ad
          14766 => x"84", -- $039ae
          14767 => x"85", -- $039af
          14768 => x"86", -- $039b0
          14769 => x"87", -- $039b1
          14770 => x"88", -- $039b2
          14771 => x"87", -- $039b3
          14772 => x"88", -- $039b4
          14773 => x"88", -- $039b5
          14774 => x"87", -- $039b6
          14775 => x"87", -- $039b7
          14776 => x"86", -- $039b8
          14777 => x"85", -- $039b9
          14778 => x"84", -- $039ba
          14779 => x"83", -- $039bb
          14780 => x"82", -- $039bc
          14781 => x"80", -- $039bd
          14782 => x"7f", -- $039be
          14783 => x"7d", -- $039bf
          14784 => x"7b", -- $039c0
          14785 => x"79", -- $039c1
          14786 => x"78", -- $039c2
          14787 => x"77", -- $039c3
          14788 => x"76", -- $039c4
          14789 => x"75", -- $039c5
          14790 => x"75", -- $039c6
          14791 => x"75", -- $039c7
          14792 => x"75", -- $039c8
          14793 => x"76", -- $039c9
          14794 => x"77", -- $039ca
          14795 => x"77", -- $039cb
          14796 => x"79", -- $039cc
          14797 => x"7b", -- $039cd
          14798 => x"7c", -- $039ce
          14799 => x"7e", -- $039cf
          14800 => x"80", -- $039d0
          14801 => x"81", -- $039d1
          14802 => x"82", -- $039d2
          14803 => x"83", -- $039d3
          14804 => x"85", -- $039d4
          14805 => x"86", -- $039d5
          14806 => x"87", -- $039d6
          14807 => x"88", -- $039d7
          14808 => x"88", -- $039d8
          14809 => x"89", -- $039d9
          14810 => x"89", -- $039da
          14811 => x"8a", -- $039db
          14812 => x"8a", -- $039dc
          14813 => x"89", -- $039dd
          14814 => x"8a", -- $039de
          14815 => x"89", -- $039df
          14816 => x"88", -- $039e0
          14817 => x"87", -- $039e1
          14818 => x"86", -- $039e2
          14819 => x"85", -- $039e3
          14820 => x"83", -- $039e4
          14821 => x"82", -- $039e5
          14822 => x"81", -- $039e6
          14823 => x"7f", -- $039e7
          14824 => x"7c", -- $039e8
          14825 => x"7b", -- $039e9
          14826 => x"78", -- $039ea
          14827 => x"76", -- $039eb
          14828 => x"74", -- $039ec
          14829 => x"73", -- $039ed
          14830 => x"72", -- $039ee
          14831 => x"71", -- $039ef
          14832 => x"71", -- $039f0
          14833 => x"71", -- $039f1
          14834 => x"72", -- $039f2
          14835 => x"74", -- $039f3
          14836 => x"76", -- $039f4
          14837 => x"78", -- $039f5
          14838 => x"7a", -- $039f6
          14839 => x"7e", -- $039f7
          14840 => x"80", -- $039f8
          14841 => x"81", -- $039f9
          14842 => x"83", -- $039fa
          14843 => x"85", -- $039fb
          14844 => x"86", -- $039fc
          14845 => x"87", -- $039fd
          14846 => x"87", -- $039fe
          14847 => x"86", -- $039ff
          14848 => x"85", -- $03a00
          14849 => x"84", -- $03a01
          14850 => x"83", -- $03a02
          14851 => x"81", -- $03a03
          14852 => x"81", -- $03a04
          14853 => x"81", -- $03a05
          14854 => x"80", -- $03a06
          14855 => x"80", -- $03a07
          14856 => x"81", -- $03a08
          14857 => x"82", -- $03a09
          14858 => x"82", -- $03a0a
          14859 => x"83", -- $03a0b
          14860 => x"84", -- $03a0c
          14861 => x"84", -- $03a0d
          14862 => x"85", -- $03a0e
          14863 => x"84", -- $03a0f
          14864 => x"83", -- $03a10
          14865 => x"82", -- $03a11
          14866 => x"81", -- $03a12
          14867 => x"80", -- $03a13
          14868 => x"7e", -- $03a14
          14869 => x"7d", -- $03a15
          14870 => x"7c", -- $03a16
          14871 => x"7a", -- $03a17
          14872 => x"79", -- $03a18
          14873 => x"78", -- $03a19
          14874 => x"77", -- $03a1a
          14875 => x"77", -- $03a1b
          14876 => x"77", -- $03a1c
          14877 => x"77", -- $03a1d
          14878 => x"77", -- $03a1e
          14879 => x"77", -- $03a1f
          14880 => x"78", -- $03a20
          14881 => x"79", -- $03a21
          14882 => x"79", -- $03a22
          14883 => x"7a", -- $03a23
          14884 => x"7c", -- $03a24
          14885 => x"7c", -- $03a25
          14886 => x"7d", -- $03a26
          14887 => x"7e", -- $03a27
          14888 => x"7f", -- $03a28
          14889 => x"7f", -- $03a29
          14890 => x"80", -- $03a2a
          14891 => x"80", -- $03a2b
          14892 => x"80", -- $03a2c
          14893 => x"81", -- $03a2d
          14894 => x"83", -- $03a2e
          14895 => x"83", -- $03a2f
          14896 => x"83", -- $03a30
          14897 => x"84", -- $03a31
          14898 => x"84", -- $03a32
          14899 => x"84", -- $03a33
          14900 => x"85", -- $03a34
          14901 => x"87", -- $03a35
          14902 => x"87", -- $03a36
          14903 => x"88", -- $03a37
          14904 => x"89", -- $03a38
          14905 => x"87", -- $03a39
          14906 => x"88", -- $03a3a
          14907 => x"88", -- $03a3b
          14908 => x"84", -- $03a3c
          14909 => x"85", -- $03a3d
          14910 => x"84", -- $03a3e
          14911 => x"82", -- $03a3f
          14912 => x"80", -- $03a40
          14913 => x"80", -- $03a41
          14914 => x"7e", -- $03a42
          14915 => x"79", -- $03a43
          14916 => x"78", -- $03a44
          14917 => x"77", -- $03a45
          14918 => x"73", -- $03a46
          14919 => x"72", -- $03a47
          14920 => x"74", -- $03a48
          14921 => x"73", -- $03a49
          14922 => x"71", -- $03a4a
          14923 => x"74", -- $03a4b
          14924 => x"75", -- $03a4c
          14925 => x"76", -- $03a4d
          14926 => x"79", -- $03a4e
          14927 => x"7c", -- $03a4f
          14928 => x"7e", -- $03a50
          14929 => x"80", -- $03a51
          14930 => x"82", -- $03a52
          14931 => x"83", -- $03a53
          14932 => x"85", -- $03a54
          14933 => x"86", -- $03a55
          14934 => x"87", -- $03a56
          14935 => x"87", -- $03a57
          14936 => x"86", -- $03a58
          14937 => x"85", -- $03a59
          14938 => x"83", -- $03a5a
          14939 => x"82", -- $03a5b
          14940 => x"80", -- $03a5c
          14941 => x"7f", -- $03a5d
          14942 => x"7e", -- $03a5e
          14943 => x"7c", -- $03a5f
          14944 => x"7c", -- $03a60
          14945 => x"7b", -- $03a61
          14946 => x"7c", -- $03a62
          14947 => x"7c", -- $03a63
          14948 => x"7e", -- $03a64
          14949 => x"7f", -- $03a65
          14950 => x"80", -- $03a66
          14951 => x"80", -- $03a67
          14952 => x"82", -- $03a68
          14953 => x"83", -- $03a69
          14954 => x"82", -- $03a6a
          14955 => x"83", -- $03a6b
          14956 => x"83", -- $03a6c
          14957 => x"82", -- $03a6d
          14958 => x"81", -- $03a6e
          14959 => x"81", -- $03a6f
          14960 => x"80", -- $03a70
          14961 => x"80", -- $03a71
          14962 => x"80", -- $03a72
          14963 => x"80", -- $03a73
          14964 => x"80", -- $03a74
          14965 => x"80", -- $03a75
          14966 => x"80", -- $03a76
          14967 => x"80", -- $03a77
          14968 => x"80", -- $03a78
          14969 => x"80", -- $03a79
          14970 => x"7f", -- $03a7a
          14971 => x"7f", -- $03a7b
          14972 => x"7f", -- $03a7c
          14973 => x"7d", -- $03a7d
          14974 => x"7d", -- $03a7e
          14975 => x"7d", -- $03a7f
          14976 => x"7b", -- $03a80
          14977 => x"7a", -- $03a81
          14978 => x"7a", -- $03a82
          14979 => x"79", -- $03a83
          14980 => x"78", -- $03a84
          14981 => x"79", -- $03a85
          14982 => x"79", -- $03a86
          14983 => x"78", -- $03a87
          14984 => x"78", -- $03a88
          14985 => x"7a", -- $03a89
          14986 => x"7a", -- $03a8a
          14987 => x"7a", -- $03a8b
          14988 => x"7d", -- $03a8c
          14989 => x"7e", -- $03a8d
          14990 => x"7f", -- $03a8e
          14991 => x"80", -- $03a8f
          14992 => x"81", -- $03a90
          14993 => x"82", -- $03a91
          14994 => x"84", -- $03a92
          14995 => x"86", -- $03a93
          14996 => x"88", -- $03a94
          14997 => x"89", -- $03a95
          14998 => x"8b", -- $03a96
          14999 => x"8a", -- $03a97
          15000 => x"8a", -- $03a98
          15001 => x"89", -- $03a99
          15002 => x"87", -- $03a9a
          15003 => x"87", -- $03a9b
          15004 => x"86", -- $03a9c
          15005 => x"84", -- $03a9d
          15006 => x"82", -- $03a9e
          15007 => x"81", -- $03a9f
          15008 => x"80", -- $03aa0
          15009 => x"7c", -- $03aa1
          15010 => x"7c", -- $03aa2
          15011 => x"7b", -- $03aa3
          15012 => x"79", -- $03aa4
          15013 => x"78", -- $03aa5
          15014 => x"78", -- $03aa6
          15015 => x"78", -- $03aa7
          15016 => x"77", -- $03aa8
          15017 => x"78", -- $03aa9
          15018 => x"78", -- $03aaa
          15019 => x"78", -- $03aab
          15020 => x"79", -- $03aac
          15021 => x"7a", -- $03aad
          15022 => x"7b", -- $03aae
          15023 => x"7c", -- $03aaf
          15024 => x"7d", -- $03ab0
          15025 => x"7e", -- $03ab1
          15026 => x"7f", -- $03ab2
          15027 => x"80", -- $03ab3
          15028 => x"80", -- $03ab4
          15029 => x"80", -- $03ab5
          15030 => x"80", -- $03ab6
          15031 => x"80", -- $03ab7
          15032 => x"80", -- $03ab8
          15033 => x"7f", -- $03ab9
          15034 => x"7e", -- $03aba
          15035 => x"7d", -- $03abb
          15036 => x"7d", -- $03abc
          15037 => x"7c", -- $03abd
          15038 => x"7c", -- $03abe
          15039 => x"7c", -- $03abf
          15040 => x"7d", -- $03ac0
          15041 => x"7e", -- $03ac1
          15042 => x"7f", -- $03ac2
          15043 => x"80", -- $03ac3
          15044 => x"81", -- $03ac4
          15045 => x"83", -- $03ac5
          15046 => x"84", -- $03ac6
          15047 => x"84", -- $03ac7
          15048 => x"85", -- $03ac8
          15049 => x"85", -- $03ac9
          15050 => x"86", -- $03aca
          15051 => x"86", -- $03acb
          15052 => x"85", -- $03acc
          15053 => x"85", -- $03acd
          15054 => x"84", -- $03ace
          15055 => x"83", -- $03acf
          15056 => x"82", -- $03ad0
          15057 => x"82", -- $03ad1
          15058 => x"81", -- $03ad2
          15059 => x"80", -- $03ad3
          15060 => x"80", -- $03ad4
          15061 => x"80", -- $03ad5
          15062 => x"7f", -- $03ad6
          15063 => x"7e", -- $03ad7
          15064 => x"7e", -- $03ad8
          15065 => x"7d", -- $03ad9
          15066 => x"7b", -- $03ada
          15067 => x"7b", -- $03adb
          15068 => x"7a", -- $03adc
          15069 => x"78", -- $03add
          15070 => x"78", -- $03ade
          15071 => x"77", -- $03adf
          15072 => x"76", -- $03ae0
          15073 => x"75", -- $03ae1
          15074 => x"75", -- $03ae2
          15075 => x"75", -- $03ae3
          15076 => x"76", -- $03ae4
          15077 => x"76", -- $03ae5
          15078 => x"77", -- $03ae6
          15079 => x"79", -- $03ae7
          15080 => x"7b", -- $03ae8
          15081 => x"7c", -- $03ae9
          15082 => x"7e", -- $03aea
          15083 => x"80", -- $03aeb
          15084 => x"82", -- $03aec
          15085 => x"84", -- $03aed
          15086 => x"86", -- $03aee
          15087 => x"88", -- $03aef
          15088 => x"8a", -- $03af0
          15089 => x"8b", -- $03af1
          15090 => x"8c", -- $03af2
          15091 => x"8d", -- $03af3
          15092 => x"8e", -- $03af4
          15093 => x"8e", -- $03af5
          15094 => x"8d", -- $03af6
          15095 => x"8b", -- $03af7
          15096 => x"8a", -- $03af8
          15097 => x"87", -- $03af9
          15098 => x"84", -- $03afa
          15099 => x"83", -- $03afb
          15100 => x"82", -- $03afc
          15101 => x"80", -- $03afd
          15102 => x"7e", -- $03afe
          15103 => x"7e", -- $03aff
          15104 => x"7b", -- $03b00
          15105 => x"79", -- $03b01
          15106 => x"79", -- $03b02
          15107 => x"77", -- $03b03
          15108 => x"76", -- $03b04
          15109 => x"77", -- $03b05
          15110 => x"76", -- $03b06
          15111 => x"76", -- $03b07
          15112 => x"76", -- $03b08
          15113 => x"77", -- $03b09
          15114 => x"77", -- $03b0a
          15115 => x"78", -- $03b0b
          15116 => x"79", -- $03b0c
          15117 => x"7a", -- $03b0d
          15118 => x"7b", -- $03b0e
          15119 => x"7d", -- $03b0f
          15120 => x"7f", -- $03b10
          15121 => x"80", -- $03b11
          15122 => x"81", -- $03b12
          15123 => x"82", -- $03b13
          15124 => x"82", -- $03b14
          15125 => x"83", -- $03b15
          15126 => x"83", -- $03b16
          15127 => x"83", -- $03b17
          15128 => x"83", -- $03b18
          15129 => x"82", -- $03b19
          15130 => x"81", -- $03b1a
          15131 => x"81", -- $03b1b
          15132 => x"80", -- $03b1c
          15133 => x"80", -- $03b1d
          15134 => x"80", -- $03b1e
          15135 => x"7f", -- $03b1f
          15136 => x"7f", -- $03b20
          15137 => x"80", -- $03b21
          15138 => x"80", -- $03b22
          15139 => x"80", -- $03b23
          15140 => x"81", -- $03b24
          15141 => x"82", -- $03b25
          15142 => x"82", -- $03b26
          15143 => x"83", -- $03b27
          15144 => x"83", -- $03b28
          15145 => x"83", -- $03b29
          15146 => x"83", -- $03b2a
          15147 => x"83", -- $03b2b
          15148 => x"83", -- $03b2c
          15149 => x"82", -- $03b2d
          15150 => x"82", -- $03b2e
          15151 => x"82", -- $03b2f
          15152 => x"82", -- $03b30
          15153 => x"82", -- $03b31
          15154 => x"83", -- $03b32
          15155 => x"82", -- $03b33
          15156 => x"82", -- $03b34
          15157 => x"82", -- $03b35
          15158 => x"82", -- $03b36
          15159 => x"81", -- $03b37
          15160 => x"81", -- $03b38
          15161 => x"80", -- $03b39
          15162 => x"80", -- $03b3a
          15163 => x"7e", -- $03b3b
          15164 => x"7d", -- $03b3c
          15165 => x"7c", -- $03b3d
          15166 => x"7a", -- $03b3e
          15167 => x"79", -- $03b3f
          15168 => x"79", -- $03b40
          15169 => x"78", -- $03b41
          15170 => x"77", -- $03b42
          15171 => x"78", -- $03b43
          15172 => x"78", -- $03b44
          15173 => x"78", -- $03b45
          15174 => x"79", -- $03b46
          15175 => x"7b", -- $03b47
          15176 => x"7b", -- $03b48
          15177 => x"7c", -- $03b49
          15178 => x"7e", -- $03b4a
          15179 => x"7f", -- $03b4b
          15180 => x"80", -- $03b4c
          15181 => x"80", -- $03b4d
          15182 => x"81", -- $03b4e
          15183 => x"82", -- $03b4f
          15184 => x"84", -- $03b50
          15185 => x"85", -- $03b51
          15186 => x"86", -- $03b52
          15187 => x"87", -- $03b53
          15188 => x"88", -- $03b54
          15189 => x"8a", -- $03b55
          15190 => x"8b", -- $03b56
          15191 => x"8c", -- $03b57
          15192 => x"8b", -- $03b58
          15193 => x"8a", -- $03b59
          15194 => x"8b", -- $03b5a
          15195 => x"88", -- $03b5b
          15196 => x"88", -- $03b5c
          15197 => x"88", -- $03b5d
          15198 => x"86", -- $03b5e
          15199 => x"85", -- $03b5f
          15200 => x"84", -- $03b60
          15201 => x"83", -- $03b61
          15202 => x"80", -- $03b62
          15203 => x"80", -- $03b63
          15204 => x"80", -- $03b64
          15205 => x"7d", -- $03b65
          15206 => x"7d", -- $03b66
          15207 => x"7c", -- $03b67
          15208 => x"7a", -- $03b68
          15209 => x"7a", -- $03b69
          15210 => x"79", -- $03b6a
          15211 => x"78", -- $03b6b
          15212 => x"78", -- $03b6c
          15213 => x"77", -- $03b6d
          15214 => x"77", -- $03b6e
          15215 => x"78", -- $03b6f
          15216 => x"79", -- $03b70
          15217 => x"7a", -- $03b71
          15218 => x"7c", -- $03b72
          15219 => x"7e", -- $03b73
          15220 => x"7f", -- $03b74
          15221 => x"80", -- $03b75
          15222 => x"82", -- $03b76
          15223 => x"82", -- $03b77
          15224 => x"82", -- $03b78
          15225 => x"83", -- $03b79
          15226 => x"82", -- $03b7a
          15227 => x"82", -- $03b7b
          15228 => x"82", -- $03b7c
          15229 => x"81", -- $03b7d
          15230 => x"80", -- $03b7e
          15231 => x"80", -- $03b7f
          15232 => x"80", -- $03b80
          15233 => x"80", -- $03b81
          15234 => x"80", -- $03b82
          15235 => x"81", -- $03b83
          15236 => x"82", -- $03b84
          15237 => x"83", -- $03b85
          15238 => x"84", -- $03b86
          15239 => x"85", -- $03b87
          15240 => x"86", -- $03b88
          15241 => x"87", -- $03b89
          15242 => x"87", -- $03b8a
          15243 => x"87", -- $03b8b
          15244 => x"86", -- $03b8c
          15245 => x"86", -- $03b8d
          15246 => x"86", -- $03b8e
          15247 => x"85", -- $03b8f
          15248 => x"84", -- $03b90
          15249 => x"84", -- $03b91
          15250 => x"83", -- $03b92
          15251 => x"82", -- $03b93
          15252 => x"82", -- $03b94
          15253 => x"81", -- $03b95
          15254 => x"81", -- $03b96
          15255 => x"80", -- $03b97
          15256 => x"80", -- $03b98
          15257 => x"80", -- $03b99
          15258 => x"80", -- $03b9a
          15259 => x"7f", -- $03b9b
          15260 => x"7e", -- $03b9c
          15261 => x"7d", -- $03b9d
          15262 => x"7c", -- $03b9e
          15263 => x"7b", -- $03b9f
          15264 => x"7a", -- $03ba0
          15265 => x"79", -- $03ba1
          15266 => x"78", -- $03ba2
          15267 => x"77", -- $03ba3
          15268 => x"77", -- $03ba4
          15269 => x"77", -- $03ba5
          15270 => x"78", -- $03ba6
          15271 => x"79", -- $03ba7
          15272 => x"7a", -- $03ba8
          15273 => x"7c", -- $03ba9
          15274 => x"7d", -- $03baa
          15275 => x"7f", -- $03bab
          15276 => x"80", -- $03bac
          15277 => x"81", -- $03bad
          15278 => x"83", -- $03bae
          15279 => x"84", -- $03baf
          15280 => x"86", -- $03bb0
          15281 => x"88", -- $03bb1
          15282 => x"89", -- $03bb2
          15283 => x"8a", -- $03bb3
          15284 => x"8b", -- $03bb4
          15285 => x"8c", -- $03bb5
          15286 => x"8d", -- $03bb6
          15287 => x"8d", -- $03bb7
          15288 => x"8d", -- $03bb8
          15289 => x"8c", -- $03bb9
          15290 => x"8b", -- $03bba
          15291 => x"8a", -- $03bbb
          15292 => x"88", -- $03bbc
          15293 => x"86", -- $03bbd
          15294 => x"84", -- $03bbe
          15295 => x"82", -- $03bbf
          15296 => x"81", -- $03bc0
          15297 => x"80", -- $03bc1
          15298 => x"7f", -- $03bc2
          15299 => x"7e", -- $03bc3
          15300 => x"7c", -- $03bc4
          15301 => x"7b", -- $03bc5
          15302 => x"7a", -- $03bc6
          15303 => x"7a", -- $03bc7
          15304 => x"7a", -- $03bc8
          15305 => x"79", -- $03bc9
          15306 => x"79", -- $03bca
          15307 => x"79", -- $03bcb
          15308 => x"78", -- $03bcc
          15309 => x"78", -- $03bcd
          15310 => x"78", -- $03bce
          15311 => x"79", -- $03bcf
          15312 => x"7a", -- $03bd0
          15313 => x"7a", -- $03bd1
          15314 => x"7b", -- $03bd2
          15315 => x"7c", -- $03bd3
          15316 => x"7d", -- $03bd4
          15317 => x"7e", -- $03bd5
          15318 => x"80", -- $03bd6
          15319 => x"80", -- $03bd7
          15320 => x"81", -- $03bd8
          15321 => x"82", -- $03bd9
          15322 => x"82", -- $03bda
          15323 => x"83", -- $03bdb
          15324 => x"83", -- $03bdc
          15325 => x"83", -- $03bdd
          15326 => x"83", -- $03bde
          15327 => x"83", -- $03bdf
          15328 => x"82", -- $03be0
          15329 => x"82", -- $03be1
          15330 => x"81", -- $03be2
          15331 => x"82", -- $03be3
          15332 => x"82", -- $03be4
          15333 => x"82", -- $03be5
          15334 => x"83", -- $03be6
          15335 => x"84", -- $03be7
          15336 => x"85", -- $03be8
          15337 => x"86", -- $03be9
          15338 => x"86", -- $03bea
          15339 => x"88", -- $03beb
          15340 => x"88", -- $03bec
          15341 => x"87", -- $03bed
          15342 => x"87", -- $03bee
          15343 => x"87", -- $03bef
          15344 => x"86", -- $03bf0
          15345 => x"85", -- $03bf1
          15346 => x"85", -- $03bf2
          15347 => x"84", -- $03bf3
          15348 => x"83", -- $03bf4
          15349 => x"83", -- $03bf5
          15350 => x"82", -- $03bf6
          15351 => x"80", -- $03bf7
          15352 => x"80", -- $03bf8
          15353 => x"80", -- $03bf9
          15354 => x"7e", -- $03bfa
          15355 => x"7e", -- $03bfb
          15356 => x"7d", -- $03bfc
          15357 => x"7b", -- $03bfd
          15358 => x"7a", -- $03bfe
          15359 => x"79", -- $03bff
          15360 => x"78", -- $03c00
          15361 => x"78", -- $03c01
          15362 => x"78", -- $03c02
          15363 => x"78", -- $03c03
          15364 => x"79", -- $03c04
          15365 => x"7a", -- $03c05
          15366 => x"7b", -- $03c06
          15367 => x"7c", -- $03c07
          15368 => x"7e", -- $03c08
          15369 => x"7f", -- $03c09
          15370 => x"80", -- $03c0a
          15371 => x"81", -- $03c0b
          15372 => x"81", -- $03c0c
          15373 => x"82", -- $03c0d
          15374 => x"83", -- $03c0e
          15375 => x"83", -- $03c0f
          15376 => x"83", -- $03c10
          15377 => x"83", -- $03c11
          15378 => x"83", -- $03c12
          15379 => x"83", -- $03c13
          15380 => x"83", -- $03c14
          15381 => x"83", -- $03c15
          15382 => x"84", -- $03c16
          15383 => x"85", -- $03c17
          15384 => x"85", -- $03c18
          15385 => x"86", -- $03c19
          15386 => x"86", -- $03c1a
          15387 => x"87", -- $03c1b
          15388 => x"86", -- $03c1c
          15389 => x"87", -- $03c1d
          15390 => x"86", -- $03c1e
          15391 => x"86", -- $03c1f
          15392 => x"85", -- $03c20
          15393 => x"84", -- $03c21
          15394 => x"84", -- $03c22
          15395 => x"83", -- $03c23
          15396 => x"82", -- $03c24
          15397 => x"81", -- $03c25
          15398 => x"81", -- $03c26
          15399 => x"81", -- $03c27
          15400 => x"81", -- $03c28
          15401 => x"81", -- $03c29
          15402 => x"82", -- $03c2a
          15403 => x"81", -- $03c2b
          15404 => x"82", -- $03c2c
          15405 => x"81", -- $03c2d
          15406 => x"80", -- $03c2e
          15407 => x"80", -- $03c2f
          15408 => x"7f", -- $03c30
          15409 => x"7e", -- $03c31
          15410 => x"7d", -- $03c32
          15411 => x"7c", -- $03c33
          15412 => x"7b", -- $03c34
          15413 => x"7a", -- $03c35
          15414 => x"79", -- $03c36
          15415 => x"78", -- $03c37
          15416 => x"78", -- $03c38
          15417 => x"78", -- $03c39
          15418 => x"79", -- $03c3a
          15419 => x"7a", -- $03c3b
          15420 => x"7b", -- $03c3c
          15421 => x"7c", -- $03c3d
          15422 => x"7e", -- $03c3e
          15423 => x"7f", -- $03c3f
          15424 => x"80", -- $03c40
          15425 => x"81", -- $03c41
          15426 => x"83", -- $03c42
          15427 => x"84", -- $03c43
          15428 => x"86", -- $03c44
          15429 => x"87", -- $03c45
          15430 => x"88", -- $03c46
          15431 => x"89", -- $03c47
          15432 => x"8b", -- $03c48
          15433 => x"8b", -- $03c49
          15434 => x"8b", -- $03c4a
          15435 => x"8c", -- $03c4b
          15436 => x"8c", -- $03c4c
          15437 => x"8c", -- $03c4d
          15438 => x"8c", -- $03c4e
          15439 => x"8a", -- $03c4f
          15440 => x"89", -- $03c50
          15441 => x"88", -- $03c51
          15442 => x"86", -- $03c52
          15443 => x"85", -- $03c53
          15444 => x"84", -- $03c54
          15445 => x"82", -- $03c55
          15446 => x"80", -- $03c56
          15447 => x"7f", -- $03c57
          15448 => x"7d", -- $03c58
          15449 => x"7b", -- $03c59
          15450 => x"7b", -- $03c5a
          15451 => x"79", -- $03c5b
          15452 => x"78", -- $03c5c
          15453 => x"78", -- $03c5d
          15454 => x"77", -- $03c5e
          15455 => x"77", -- $03c5f
          15456 => x"77", -- $03c60
          15457 => x"77", -- $03c61
          15458 => x"77", -- $03c62
          15459 => x"78", -- $03c63
          15460 => x"78", -- $03c64
          15461 => x"79", -- $03c65
          15462 => x"7a", -- $03c66
          15463 => x"7c", -- $03c67
          15464 => x"7d", -- $03c68
          15465 => x"7f", -- $03c69
          15466 => x"80", -- $03c6a
          15467 => x"81", -- $03c6b
          15468 => x"82", -- $03c6c
          15469 => x"83", -- $03c6d
          15470 => x"83", -- $03c6e
          15471 => x"84", -- $03c6f
          15472 => x"84", -- $03c70
          15473 => x"84", -- $03c71
          15474 => x"84", -- $03c72
          15475 => x"83", -- $03c73
          15476 => x"83", -- $03c74
          15477 => x"82", -- $03c75
          15478 => x"82", -- $03c76
          15479 => x"81", -- $03c77
          15480 => x"81", -- $03c78
          15481 => x"82", -- $03c79
          15482 => x"82", -- $03c7a
          15483 => x"83", -- $03c7b
          15484 => x"83", -- $03c7c
          15485 => x"84", -- $03c7d
          15486 => x"84", -- $03c7e
          15487 => x"85", -- $03c7f
          15488 => x"85", -- $03c80
          15489 => x"85", -- $03c81
          15490 => x"85", -- $03c82
          15491 => x"84", -- $03c83
          15492 => x"84", -- $03c84
          15493 => x"83", -- $03c85
          15494 => x"82", -- $03c86
          15495 => x"82", -- $03c87
          15496 => x"81", -- $03c88
          15497 => x"80", -- $03c89
          15498 => x"80", -- $03c8a
          15499 => x"80", -- $03c8b
          15500 => x"7f", -- $03c8c
          15501 => x"7e", -- $03c8d
          15502 => x"7d", -- $03c8e
          15503 => x"7d", -- $03c8f
          15504 => x"7c", -- $03c90
          15505 => x"7c", -- $03c91
          15506 => x"7b", -- $03c92
          15507 => x"7a", -- $03c93
          15508 => x"7a", -- $03c94
          15509 => x"79", -- $03c95
          15510 => x"79", -- $03c96
          15511 => x"79", -- $03c97
          15512 => x"79", -- $03c98
          15513 => x"79", -- $03c99
          15514 => x"7a", -- $03c9a
          15515 => x"7b", -- $03c9b
          15516 => x"7b", -- $03c9c
          15517 => x"7d", -- $03c9d
          15518 => x"7e", -- $03c9e
          15519 => x"7f", -- $03c9f
          15520 => x"80", -- $03ca0
          15521 => x"80", -- $03ca1
          15522 => x"81", -- $03ca2
          15523 => x"82", -- $03ca3
          15524 => x"82", -- $03ca4
          15525 => x"82", -- $03ca5
          15526 => x"82", -- $03ca6
          15527 => x"83", -- $03ca7
          15528 => x"83", -- $03ca8
          15529 => x"83", -- $03ca9
          15530 => x"83", -- $03caa
          15531 => x"84", -- $03cab
          15532 => x"84", -- $03cac
          15533 => x"85", -- $03cad
          15534 => x"85", -- $03cae
          15535 => x"85", -- $03caf
          15536 => x"85", -- $03cb0
          15537 => x"86", -- $03cb1
          15538 => x"85", -- $03cb2
          15539 => x"85", -- $03cb3
          15540 => x"85", -- $03cb4
          15541 => x"84", -- $03cb5
          15542 => x"83", -- $03cb6
          15543 => x"83", -- $03cb7
          15544 => x"82", -- $03cb8
          15545 => x"81", -- $03cb9
          15546 => x"81", -- $03cba
          15547 => x"80", -- $03cbb
          15548 => x"80", -- $03cbc
          15549 => x"80", -- $03cbd
          15550 => x"80", -- $03cbe
          15551 => x"80", -- $03cbf
          15552 => x"7f", -- $03cc0
          15553 => x"7f", -- $03cc1
          15554 => x"7e", -- $03cc2
          15555 => x"7e", -- $03cc3
          15556 => x"7d", -- $03cc4
          15557 => x"7c", -- $03cc5
          15558 => x"7b", -- $03cc6
          15559 => x"7a", -- $03cc7
          15560 => x"7a", -- $03cc8
          15561 => x"7a", -- $03cc9
          15562 => x"7a", -- $03cca
          15563 => x"7a", -- $03ccb
          15564 => x"7a", -- $03ccc
          15565 => x"7a", -- $03ccd
          15566 => x"7b", -- $03cce
          15567 => x"7c", -- $03ccf
          15568 => x"7d", -- $03cd0
          15569 => x"7e", -- $03cd1
          15570 => x"7f", -- $03cd2
          15571 => x"80", -- $03cd3
          15572 => x"80", -- $03cd4
          15573 => x"81", -- $03cd5
          15574 => x"81", -- $03cd6
          15575 => x"82", -- $03cd7
          15576 => x"82", -- $03cd8
          15577 => x"82", -- $03cd9
          15578 => x"82", -- $03cda
          15579 => x"82", -- $03cdb
          15580 => x"82", -- $03cdc
          15581 => x"83", -- $03cdd
          15582 => x"83", -- $03cde
          15583 => x"84", -- $03cdf
          15584 => x"85", -- $03ce0
          15585 => x"85", -- $03ce1
          15586 => x"86", -- $03ce2
          15587 => x"86", -- $03ce3
          15588 => x"86", -- $03ce4
          15589 => x"86", -- $03ce5
          15590 => x"86", -- $03ce6
          15591 => x"86", -- $03ce7
          15592 => x"84", -- $03ce8
          15593 => x"84", -- $03ce9
          15594 => x"83", -- $03cea
          15595 => x"81", -- $03ceb
          15596 => x"81", -- $03cec
          15597 => x"80", -- $03ced
          15598 => x"80", -- $03cee
          15599 => x"7f", -- $03cef
          15600 => x"7f", -- $03cf0
          15601 => x"7e", -- $03cf1
          15602 => x"7e", -- $03cf2
          15603 => x"7d", -- $03cf3
          15604 => x"7c", -- $03cf4
          15605 => x"7c", -- $03cf5
          15606 => x"7b", -- $03cf6
          15607 => x"7a", -- $03cf7
          15608 => x"79", -- $03cf8
          15609 => x"79", -- $03cf9
          15610 => x"78", -- $03cfa
          15611 => x"78", -- $03cfb
          15612 => x"78", -- $03cfc
          15613 => x"78", -- $03cfd
          15614 => x"78", -- $03cfe
          15615 => x"79", -- $03cff
          15616 => x"7a", -- $03d00
          15617 => x"7b", -- $03d01
          15618 => x"7d", -- $03d02
          15619 => x"7e", -- $03d03
          15620 => x"7f", -- $03d04
          15621 => x"80", -- $03d05
          15622 => x"81", -- $03d06
          15623 => x"81", -- $03d07
          15624 => x"82", -- $03d08
          15625 => x"82", -- $03d09
          15626 => x"83", -- $03d0a
          15627 => x"82", -- $03d0b
          15628 => x"82", -- $03d0c
          15629 => x"82", -- $03d0d
          15630 => x"82", -- $03d0e
          15631 => x"82", -- $03d0f
          15632 => x"83", -- $03d10
          15633 => x"83", -- $03d11
          15634 => x"84", -- $03d12
          15635 => x"84", -- $03d13
          15636 => x"85", -- $03d14
          15637 => x"85", -- $03d15
          15638 => x"86", -- $03d16
          15639 => x"86", -- $03d17
          15640 => x"86", -- $03d18
          15641 => x"85", -- $03d19
          15642 => x"84", -- $03d1a
          15643 => x"83", -- $03d1b
          15644 => x"82", -- $03d1c
          15645 => x"81", -- $03d1d
          15646 => x"80", -- $03d1e
          15647 => x"80", -- $03d1f
          15648 => x"7f", -- $03d20
          15649 => x"7e", -- $03d21
          15650 => x"7d", -- $03d22
          15651 => x"7c", -- $03d23
          15652 => x"7c", -- $03d24
          15653 => x"7b", -- $03d25
          15654 => x"7b", -- $03d26
          15655 => x"7b", -- $03d27
          15656 => x"7b", -- $03d28
          15657 => x"7a", -- $03d29
          15658 => x"7a", -- $03d2a
          15659 => x"79", -- $03d2b
          15660 => x"79", -- $03d2c
          15661 => x"79", -- $03d2d
          15662 => x"79", -- $03d2e
          15663 => x"79", -- $03d2f
          15664 => x"79", -- $03d30
          15665 => x"7a", -- $03d31
          15666 => x"7b", -- $03d32
          15667 => x"7c", -- $03d33
          15668 => x"7d", -- $03d34
          15669 => x"7f", -- $03d35
          15670 => x"80", -- $03d36
          15671 => x"80", -- $03d37
          15672 => x"82", -- $03d38
          15673 => x"83", -- $03d39
          15674 => x"83", -- $03d3a
          15675 => x"83", -- $03d3b
          15676 => x"84", -- $03d3c
          15677 => x"84", -- $03d3d
          15678 => x"84", -- $03d3e
          15679 => x"83", -- $03d3f
          15680 => x"83", -- $03d40
          15681 => x"82", -- $03d41
          15682 => x"82", -- $03d42
          15683 => x"82", -- $03d43
          15684 => x"82", -- $03d44
          15685 => x"82", -- $03d45
          15686 => x"82", -- $03d46
          15687 => x"82", -- $03d47
          15688 => x"82", -- $03d48
          15689 => x"82", -- $03d49
          15690 => x"82", -- $03d4a
          15691 => x"82", -- $03d4b
          15692 => x"82", -- $03d4c
          15693 => x"81", -- $03d4d
          15694 => x"81", -- $03d4e
          15695 => x"80", -- $03d4f
          15696 => x"80", -- $03d50
          15697 => x"7f", -- $03d51
          15698 => x"7f", -- $03d52
          15699 => x"7e", -- $03d53
          15700 => x"7e", -- $03d54
          15701 => x"7e", -- $03d55
          15702 => x"7e", -- $03d56
          15703 => x"7e", -- $03d57
          15704 => x"7e", -- $03d58
          15705 => x"7e", -- $03d59
          15706 => x"7e", -- $03d5a
          15707 => x"7e", -- $03d5b
          15708 => x"7d", -- $03d5c
          15709 => x"7d", -- $03d5d
          15710 => x"7c", -- $03d5e
          15711 => x"7b", -- $03d5f
          15712 => x"7b", -- $03d60
          15713 => x"7a", -- $03d61
          15714 => x"7a", -- $03d62
          15715 => x"7a", -- $03d63
          15716 => x"7a", -- $03d64
          15717 => x"7b", -- $03d65
          15718 => x"7b", -- $03d66
          15719 => x"7c", -- $03d67
          15720 => x"7d", -- $03d68
          15721 => x"7e", -- $03d69
          15722 => x"7f", -- $03d6a
          15723 => x"80", -- $03d6b
          15724 => x"80", -- $03d6c
          15725 => x"81", -- $03d6d
          15726 => x"81", -- $03d6e
          15727 => x"82", -- $03d6f
          15728 => x"82", -- $03d70
          15729 => x"82", -- $03d71
          15730 => x"82", -- $03d72
          15731 => x"82", -- $03d73
          15732 => x"82", -- $03d74
          15733 => x"82", -- $03d75
          15734 => x"82", -- $03d76
          15735 => x"83", -- $03d77
          15736 => x"83", -- $03d78
          15737 => x"83", -- $03d79
          15738 => x"83", -- $03d7a
          15739 => x"84", -- $03d7b
          15740 => x"84", -- $03d7c
          15741 => x"84", -- $03d7d
          15742 => x"84", -- $03d7e
          15743 => x"83", -- $03d7f
          15744 => x"83", -- $03d80
          15745 => x"82", -- $03d81
          15746 => x"81", -- $03d82
          15747 => x"80", -- $03d83
          15748 => x"80", -- $03d84
          15749 => x"80", -- $03d85
          15750 => x"7f", -- $03d86
          15751 => x"7f", -- $03d87
          15752 => x"7e", -- $03d88
          15753 => x"7e", -- $03d89
          15754 => x"7d", -- $03d8a
          15755 => x"7d", -- $03d8b
          15756 => x"7c", -- $03d8c
          15757 => x"7c", -- $03d8d
          15758 => x"7b", -- $03d8e
          15759 => x"7a", -- $03d8f
          15760 => x"7a", -- $03d90
          15761 => x"79", -- $03d91
          15762 => x"78", -- $03d92
          15763 => x"78", -- $03d93
          15764 => x"78", -- $03d94
          15765 => x"77", -- $03d95
          15766 => x"78", -- $03d96
          15767 => x"78", -- $03d97
          15768 => x"79", -- $03d98
          15769 => x"7b", -- $03d99
          15770 => x"7c", -- $03d9a
          15771 => x"7d", -- $03d9b
          15772 => x"7f", -- $03d9c
          15773 => x"80", -- $03d9d
          15774 => x"80", -- $03d9e
          15775 => x"81", -- $03d9f
          15776 => x"82", -- $03da0
          15777 => x"83", -- $03da1
          15778 => x"84", -- $03da2
          15779 => x"85", -- $03da3
          15780 => x"85", -- $03da4
          15781 => x"85", -- $03da5
          15782 => x"85", -- $03da6
          15783 => x"85", -- $03da7
          15784 => x"85", -- $03da8
          15785 => x"85", -- $03da9
          15786 => x"85", -- $03daa
          15787 => x"85", -- $03dab
          15788 => x"85", -- $03dac
          15789 => x"84", -- $03dad
          15790 => x"84", -- $03dae
          15791 => x"84", -- $03daf
          15792 => x"83", -- $03db0
          15793 => x"82", -- $03db1
          15794 => x"81", -- $03db2
          15795 => x"80", -- $03db3
          15796 => x"80", -- $03db4
          15797 => x"7f", -- $03db5
          15798 => x"7e", -- $03db6
          15799 => x"7e", -- $03db7
          15800 => x"7d", -- $03db8
          15801 => x"7c", -- $03db9
          15802 => x"7c", -- $03dba
          15803 => x"7b", -- $03dbb
          15804 => x"7b", -- $03dbc
          15805 => x"7b", -- $03dbd
          15806 => x"7b", -- $03dbe
          15807 => x"7b", -- $03dbf
          15808 => x"7b", -- $03dc0
          15809 => x"7b", -- $03dc1
          15810 => x"7b", -- $03dc2
          15811 => x"7b", -- $03dc3
          15812 => x"7b", -- $03dc4
          15813 => x"7b", -- $03dc5
          15814 => x"7b", -- $03dc6
          15815 => x"7b", -- $03dc7
          15816 => x"7b", -- $03dc8
          15817 => x"7c", -- $03dc9
          15818 => x"7c", -- $03dca
          15819 => x"7d", -- $03dcb
          15820 => x"7e", -- $03dcc
          15821 => x"7f", -- $03dcd
          15822 => x"80", -- $03dce
          15823 => x"81", -- $03dcf
          15824 => x"82", -- $03dd0
          15825 => x"83", -- $03dd1
          15826 => x"83", -- $03dd2
          15827 => x"84", -- $03dd3
          15828 => x"84", -- $03dd4
          15829 => x"85", -- $03dd5
          15830 => x"85", -- $03dd6
          15831 => x"85", -- $03dd7
          15832 => x"85", -- $03dd8
          15833 => x"84", -- $03dd9
          15834 => x"84", -- $03dda
          15835 => x"84", -- $03ddb
          15836 => x"83", -- $03ddc
          15837 => x"83", -- $03ddd
          15838 => x"83", -- $03dde
          15839 => x"83", -- $03ddf
          15840 => x"82", -- $03de0
          15841 => x"82", -- $03de1
          15842 => x"82", -- $03de2
          15843 => x"81", -- $03de3
          15844 => x"81", -- $03de4
          15845 => x"80", -- $03de5
          15846 => x"80", -- $03de6
          15847 => x"80", -- $03de7
          15848 => x"7f", -- $03de8
          15849 => x"7e", -- $03de9
          15850 => x"7e", -- $03dea
          15851 => x"7d", -- $03deb
          15852 => x"7d", -- $03dec
          15853 => x"7d", -- $03ded
          15854 => x"7c", -- $03dee
          15855 => x"7c", -- $03def
          15856 => x"7c", -- $03df0
          15857 => x"7c", -- $03df1
          15858 => x"7c", -- $03df2
          15859 => x"7d", -- $03df3
          15860 => x"7d", -- $03df4
          15861 => x"7d", -- $03df5
          15862 => x"7d", -- $03df6
          15863 => x"7d", -- $03df7
          15864 => x"7d", -- $03df8
          15865 => x"7d", -- $03df9
          15866 => x"7d", -- $03dfa
          15867 => x"7d", -- $03dfb
          15868 => x"7e", -- $03dfc
          15869 => x"7e", -- $03dfd
          15870 => x"7f", -- $03dfe
          15871 => x"80", -- $03dff
          15872 => x"80", -- $03e00
          15873 => x"80", -- $03e01
          15874 => x"81", -- $03e02
          15875 => x"81", -- $03e03
          15876 => x"82", -- $03e04
          15877 => x"82", -- $03e05
          15878 => x"83", -- $03e06
          15879 => x"83", -- $03e07
          15880 => x"83", -- $03e08
          15881 => x"84", -- $03e09
          15882 => x"84", -- $03e0a
          15883 => x"84", -- $03e0b
          15884 => x"84", -- $03e0c
          15885 => x"83", -- $03e0d
          15886 => x"83", -- $03e0e
          15887 => x"83", -- $03e0f
          15888 => x"83", -- $03e10
          15889 => x"83", -- $03e11
          15890 => x"82", -- $03e12
          15891 => x"82", -- $03e13
          15892 => x"81", -- $03e14
          15893 => x"81", -- $03e15
          15894 => x"80", -- $03e16
          15895 => x"80", -- $03e17
          15896 => x"80", -- $03e18
          15897 => x"80", -- $03e19
          15898 => x"7f", -- $03e1a
          15899 => x"7f", -- $03e1b
          15900 => x"7e", -- $03e1c
          15901 => x"7e", -- $03e1d
          15902 => x"7e", -- $03e1e
          15903 => x"7d", -- $03e1f
          15904 => x"7d", -- $03e20
          15905 => x"7d", -- $03e21
          15906 => x"7d", -- $03e22
          15907 => x"7d", -- $03e23
          15908 => x"7d", -- $03e24
          15909 => x"7d", -- $03e25
          15910 => x"7e", -- $03e26
          15911 => x"7d", -- $03e27
          15912 => x"7d", -- $03e28
          15913 => x"7d", -- $03e29
          15914 => x"7d", -- $03e2a
          15915 => x"7d", -- $03e2b
          15916 => x"7d", -- $03e2c
          15917 => x"7e", -- $03e2d
          15918 => x"7e", -- $03e2e
          15919 => x"7e", -- $03e2f
          15920 => x"7e", -- $03e30
          15921 => x"7f", -- $03e31
          15922 => x"7f", -- $03e32
          15923 => x"80", -- $03e33
          15924 => x"80", -- $03e34
          15925 => x"80", -- $03e35
          15926 => x"81", -- $03e36
          15927 => x"82", -- $03e37
          15928 => x"82", -- $03e38
          15929 => x"83", -- $03e39
          15930 => x"83", -- $03e3a
          15931 => x"83", -- $03e3b
          15932 => x"84", -- $03e3c
          15933 => x"84", -- $03e3d
          15934 => x"84", -- $03e3e
          15935 => x"84", -- $03e3f
          15936 => x"84", -- $03e40
          15937 => x"84", -- $03e41
          15938 => x"83", -- $03e42
          15939 => x"83", -- $03e43
          15940 => x"83", -- $03e44
          15941 => x"82", -- $03e45
          15942 => x"81", -- $03e46
          15943 => x"81", -- $03e47
          15944 => x"80", -- $03e48
          15945 => x"80", -- $03e49
          15946 => x"80", -- $03e4a
          15947 => x"7f", -- $03e4b
          15948 => x"7f", -- $03e4c
          15949 => x"7e", -- $03e4d
          15950 => x"7e", -- $03e4e
          15951 => x"7e", -- $03e4f
          15952 => x"7e", -- $03e50
          15953 => x"7d", -- $03e51
          15954 => x"7d", -- $03e52
          15955 => x"7d", -- $03e53
          15956 => x"7d", -- $03e54
          15957 => x"7d", -- $03e55
          15958 => x"7d", -- $03e56
          15959 => x"7d", -- $03e57
          15960 => x"7e", -- $03e58
          15961 => x"7e", -- $03e59
          15962 => x"7e", -- $03e5a
          15963 => x"7e", -- $03e5b
          15964 => x"7f", -- $03e5c
          15965 => x"7f", -- $03e5d
          15966 => x"7f", -- $03e5e
          15967 => x"7f", -- $03e5f
          15968 => x"7f", -- $03e60
          15969 => x"80", -- $03e61
          15970 => x"80", -- $03e62
          15971 => x"80", -- $03e63
          15972 => x"80", -- $03e64
          15973 => x"80", -- $03e65
          15974 => x"80", -- $03e66
          15975 => x"81", -- $03e67
          15976 => x"81", -- $03e68
          15977 => x"82", -- $03e69
          15978 => x"83", -- $03e6a
          15979 => x"83", -- $03e6b
          15980 => x"84", -- $03e6c
          15981 => x"84", -- $03e6d
          15982 => x"85", -- $03e6e
          15983 => x"85", -- $03e6f
          15984 => x"85", -- $03e70
          15985 => x"85", -- $03e71
          15986 => x"84", -- $03e72
          15987 => x"84", -- $03e73
          15988 => x"84", -- $03e74
          15989 => x"83", -- $03e75
          15990 => x"83", -- $03e76
          15991 => x"82", -- $03e77
          15992 => x"81", -- $03e78
          15993 => x"81", -- $03e79
          15994 => x"80", -- $03e7a
          15995 => x"80", -- $03e7b
          15996 => x"80", -- $03e7c
          15997 => x"80", -- $03e7d
          15998 => x"7f", -- $03e7e
          15999 => x"7f", -- $03e7f
          16000 => x"7f", -- $03e80
          16001 => x"7f", -- $03e81
          16002 => x"7f", -- $03e82
          16003 => x"7f", -- $03e83
          16004 => x"7f", -- $03e84
          16005 => x"7f", -- $03e85
          16006 => x"7f", -- $03e86
          16007 => x"7f", -- $03e87
          16008 => x"80", -- $03e88
          16009 => x"80", -- $03e89
          16010 => x"80", -- $03e8a
          16011 => x"80", -- $03e8b
          16012 => x"80", -- $03e8c
          16013 => x"80", -- $03e8d
          16014 => x"80", -- $03e8e
          16015 => x"80", -- $03e8f
          16016 => x"81", -- $03e90
          16017 => x"81", -- $03e91
          16018 => x"81", -- $03e92
          16019 => x"81", -- $03e93
          16020 => x"81", -- $03e94
          16021 => x"82", -- $03e95
          16022 => x"82", -- $03e96
          16023 => x"82", -- $03e97
          16024 => x"82", -- $03e98
          16025 => x"82", -- $03e99
          16026 => x"82", -- $03e9a
          16027 => x"82", -- $03e9b
          16028 => x"82", -- $03e9c
          16029 => x"82", -- $03e9d
          16030 => x"83", -- $03e9e
          16031 => x"83", -- $03e9f
          16032 => x"83", -- $03ea0
          16033 => x"83", -- $03ea1
          16034 => x"83", -- $03ea2
          16035 => x"82", -- $03ea3
          16036 => x"82", -- $03ea4
          16037 => x"82", -- $03ea5
          16038 => x"82", -- $03ea6
          16039 => x"82", -- $03ea7
          16040 => x"81", -- $03ea8
          16041 => x"81", -- $03ea9
          16042 => x"81", -- $03eaa
          16043 => x"81", -- $03eab
          16044 => x"80", -- $03eac
          16045 => x"80", -- $03ead
          16046 => x"80", -- $03eae
          16047 => x"80", -- $03eaf
          16048 => x"80", -- $03eb0
          16049 => x"80", -- $03eb1
          16050 => x"80", -- $03eb2
          16051 => x"80", -- $03eb3
          16052 => x"80", -- $03eb4
          16053 => x"80", -- $03eb5
          16054 => x"80", -- $03eb6
          16055 => x"80", -- $03eb7
          16056 => x"80", -- $03eb8
          16057 => x"80", -- $03eb9
          16058 => x"80", -- $03eba
          16059 => x"80", -- $03ebb
          16060 => x"80", -- $03ebc
          16061 => x"80", -- $03ebd
          16062 => x"80", -- $03ebe
          16063 => x"80", -- $03ebf
          16064 => x"80", -- $03ec0
          16065 => x"81", -- $03ec1
          16066 => x"81", -- $03ec2
          16067 => x"80", -- $03ec3
          16068 => x"80", -- $03ec4
          16069 => x"80", -- $03ec5
          16070 => x"80", -- $03ec6
          16071 => x"80", -- $03ec7
          16072 => x"80", -- $03ec8
          16073 => x"80", -- $03ec9
          16074 => x"80", -- $03eca
          16075 => x"80", -- $03ecb
          16076 => x"81", -- $03ecc
          16077 => x"81", -- $03ecd
          16078 => x"81", -- $03ece
          16079 => x"81", -- $03ecf
          16080 => x"81", -- $03ed0
          16081 => x"81", -- $03ed1
          16082 => x"81", -- $03ed2
          16083 => x"82", -- $03ed3
          16084 => x"82", -- $03ed4
          16085 => x"82", -- $03ed5
          16086 => x"82", -- $03ed6
          16087 => x"82", -- $03ed7
          16088 => x"82", -- $03ed8
          16089 => x"81", -- $03ed9
          16090 => x"81", -- $03eda
          16091 => x"81", -- $03edb
          16092 => x"81", -- $03edc
          16093 => x"81", -- $03edd
          16094 => x"81", -- $03ede
          16095 => x"81", -- $03edf
          16096 => x"80", -- $03ee0
          16097 => x"80", -- $03ee1
          16098 => x"80", -- $03ee2
          16099 => x"80", -- $03ee3
          16100 => x"80", -- $03ee4
          16101 => x"80", -- $03ee5
          16102 => x"80", -- $03ee6
          16103 => x"80", -- $03ee7
          16104 => x"80", -- $03ee8
          16105 => x"80", -- $03ee9
          16106 => x"80", -- $03eea
          16107 => x"80", -- $03eeb
          16108 => x"80", -- $03eec
          16109 => x"80", -- $03eed
          16110 => x"80", -- $03eee
          16111 => x"80", -- $03eef
          16112 => x"80", -- $03ef0
          16113 => x"80", -- $03ef1
          16114 => x"80", -- $03ef2
          16115 => x"80", -- $03ef3
          16116 => x"80", -- $03ef4
          16117 => x"80", -- $03ef5
          16118 => x"80", -- $03ef6
          16119 => x"80", -- $03ef7
          16120 => x"80", -- $03ef8
          16121 => x"80", -- $03ef9
          16122 => x"80", -- $03efa
          16123 => x"80", -- $03efb
          16124 => x"81", -- $03efc
          16125 => x"81", -- $03efd
          16126 => x"81", -- $03efe
          16127 => x"81", -- $03eff
          16128 => x"81", -- $03f00
          16129 => x"81", -- $03f01
          16130 => x"82", -- $03f02
          16131 => x"82", -- $03f03
          16132 => x"82", -- $03f04
          16133 => x"82", -- $03f05
          16134 => x"82", -- $03f06
          16135 => x"82", -- $03f07
          16136 => x"82", -- $03f08
          16137 => x"82", -- $03f09
          16138 => x"82", -- $03f0a
          16139 => x"82", -- $03f0b
          16140 => x"82", -- $03f0c
          16141 => x"82", -- $03f0d
          16142 => x"81", -- $03f0e
          16143 => x"81", -- $03f0f
          16144 => x"81", -- $03f10
          16145 => x"81", -- $03f11
          16146 => x"80", -- $03f12
          16147 => x"80", -- $03f13
          16148 => x"80", -- $03f14
          16149 => x"80", -- $03f15
          16150 => x"80", -- $03f16
          16151 => x"80", -- $03f17
          16152 => x"80", -- $03f18
          16153 => x"80", -- $03f19
          16154 => x"7f", -- $03f1a
          16155 => x"7f", -- $03f1b
          16156 => x"80", -- $03f1c
          16157 => x"80", -- $03f1d
          16158 => x"80", -- $03f1e
          16159 => x"80", -- $03f1f
          16160 => x"80", -- $03f20
          16161 => x"80", -- $03f21
          16162 => x"80", -- $03f22
          16163 => x"80", -- $03f23
          16164 => x"80", -- $03f24
          16165 => x"81", -- $03f25
          16166 => x"81", -- $03f26
          16167 => x"81", -- $03f27
          16168 => x"81", -- $03f28
          16169 => x"81", -- $03f29
          16170 => x"81", -- $03f2a
          16171 => x"82", -- $03f2b
          16172 => x"82", -- $03f2c
          16173 => x"82", -- $03f2d
          16174 => x"82", -- $03f2e
          16175 => x"82", -- $03f2f
          16176 => x"82", -- $03f30
          16177 => x"82", -- $03f31
          16178 => x"82", -- $03f32
          16179 => x"82", -- $03f33
          16180 => x"82", -- $03f34
          16181 => x"82", -- $03f35
          16182 => x"82", -- $03f36
          16183 => x"82", -- $03f37
          16184 => x"81", -- $03f38
          16185 => x"81", -- $03f39
          16186 => x"81", -- $03f3a
          16187 => x"81", -- $03f3b
          16188 => x"81", -- $03f3c
          16189 => x"81", -- $03f3d
          16190 => x"81", -- $03f3e
          16191 => x"81", -- $03f3f
          16192 => x"81", -- $03f40
          16193 => x"81", -- $03f41
          16194 => x"81", -- $03f42
          16195 => x"80", -- $03f43
          16196 => x"80", -- $03f44
          16197 => x"80", -- $03f45
          16198 => x"80", -- $03f46
          16199 => x"80", -- $03f47
          16200 => x"80", -- $03f48
          16201 => x"80", -- $03f49
          16202 => x"80", -- $03f4a
          16203 => x"80", -- $03f4b
          16204 => x"80", -- $03f4c
          16205 => x"80", -- $03f4d
          16206 => x"80", -- $03f4e
          16207 => x"80", -- $03f4f
          16208 => x"80", -- $03f50
          16209 => x"80", -- $03f51
          16210 => x"80", -- $03f52
          16211 => x"81", -- $03f53
          16212 => x"81", -- $03f54
          16213 => x"81", -- $03f55
          16214 => x"81", -- $03f56
          16215 => x"81", -- $03f57
          16216 => x"81", -- $03f58
          16217 => x"81", -- $03f59
          16218 => x"81", -- $03f5a
          16219 => x"81", -- $03f5b
          16220 => x"81", -- $03f5c
          16221 => x"81", -- $03f5d
          16222 => x"81", -- $03f5e
          16223 => x"81", -- $03f5f
          16224 => x"81", -- $03f60
          16225 => x"81", -- $03f61
          16226 => x"81", -- $03f62
          16227 => x"81", -- $03f63
          16228 => x"81", -- $03f64
          16229 => x"81", -- $03f65
          16230 => x"81", -- $03f66
          16231 => x"81", -- $03f67
          16232 => x"81", -- $03f68
          16233 => x"81", -- $03f69
          16234 => x"81", -- $03f6a
          16235 => x"81", -- $03f6b
          16236 => x"81", -- $03f6c
          16237 => x"81", -- $03f6d
          16238 => x"81", -- $03f6e
          16239 => x"81", -- $03f6f
          16240 => x"81", -- $03f70
          16241 => x"81", -- $03f71
          16242 => x"81", -- $03f72
          16243 => x"81", -- $03f73
          16244 => x"80", -- $03f74
          16245 => x"80", -- $03f75
          16246 => x"81", -- $03f76
          16247 => x"80", -- $03f77
          16248 => x"80", -- $03f78
          16249 => x"81", -- $03f79
          16250 => x"81", -- $03f7a
          16251 => x"80", -- $03f7b
          16252 => x"80", -- $03f7c
          16253 => x"80", -- $03f7d
          16254 => x"80", -- $03f7e
          16255 => x"80", -- $03f7f
          16256 => x"80", -- $03f80
          16257 => x"80", -- $03f81
          16258 => x"80", -- $03f82
          16259 => x"80", -- $03f83
          16260 => x"80", -- $03f84
          16261 => x"80", -- $03f85
          16262 => x"80", -- $03f86
          16263 => x"80", -- $03f87
          16264 => x"80", -- $03f88
          16265 => x"80", -- $03f89
          16266 => x"80", -- $03f8a
          16267 => x"80", -- $03f8b
          16268 => x"80", -- $03f8c
          16269 => x"80", -- $03f8d
          16270 => x"80", -- $03f8e
          16271 => x"80", -- $03f8f
          16272 => x"80", -- $03f90
          16273 => x"80", -- $03f91
          16274 => x"80", -- $03f92
          16275 => x"80", -- $03f93
          16276 => x"80", -- $03f94
          16277 => x"80", -- $03f95
          16278 => x"80", -- $03f96
          16279 => x"80", -- $03f97
          16280 => x"80", -- $03f98
          16281 => x"80", -- $03f99
          16282 => x"80", -- $03f9a
          16283 => x"80", -- $03f9b
          16284 => x"80", -- $03f9c
          16285 => x"80", -- $03f9d
          16286 => x"80", -- $03f9e
          16287 => x"80", -- $03f9f
          16288 => x"80", -- $03fa0
          16289 => x"80", -- $03fa1
          16290 => x"80", -- $03fa2
          16291 => x"80", -- $03fa3
          16292 => x"80", -- $03fa4
          16293 => x"80", -- $03fa5
          16294 => x"80", -- $03fa6
          16295 => x"80", -- $03fa7
          16296 => x"80", -- $03fa8
          16297 => x"80", -- $03fa9
          16298 => x"80", -- $03faa
          16299 => x"80", -- $03fab
          16300 => x"80", -- $03fac
          16301 => x"80", -- $03fad
          16302 => x"80", -- $03fae
          16303 => x"80", -- $03faf
          16304 => x"80", -- $03fb0
          16305 => x"80", -- $03fb1
          16306 => x"80", -- $03fb2
          16307 => x"80", -- $03fb3
          16308 => x"80", -- $03fb4
          16309 => x"80", -- $03fb5
          16310 => x"80", -- $03fb6
          16311 => x"80", -- $03fb7
          16312 => x"80", -- $03fb8
          16313 => x"80", -- $03fb9
          16314 => x"80", -- $03fba
          16315 => x"80", -- $03fbb
          16316 => x"80", -- $03fbc
          16317 => x"80", -- $03fbd
          16318 => x"80", -- $03fbe
          16319 => x"80", -- $03fbf
          16320 => x"80", -- $03fc0
          16321 => x"80", -- $03fc1
          16322 => x"80", -- $03fc2
          16323 => x"80", -- $03fc3
          16324 => x"80", -- $03fc4
          16325 => x"80", -- $03fc5
          16326 => x"80", -- $03fc6
          16327 => x"80", -- $03fc7
          16328 => x"80", -- $03fc8
          16329 => x"80", -- $03fc9
          16330 => x"80", -- $03fca
          16331 => x"80", -- $03fcb
          16332 => x"80", -- $03fcc
          16333 => x"80", -- $03fcd
          16334 => x"80", -- $03fce
          16335 => x"80", -- $03fcf
          16336 => x"80", -- $03fd0
          16337 => x"80", -- $03fd1
          16338 => x"80", -- $03fd2
          16339 => x"80", -- $03fd3
          16340 => x"80", -- $03fd4
          16341 => x"80", -- $03fd5
          16342 => x"80", -- $03fd6
          16343 => x"80", -- $03fd7
          16344 => x"80", -- $03fd8
          16345 => x"80", -- $03fd9
          16346 => x"7f", -- $03fda
          16347 => x"7f", -- $03fdb
          16348 => x"7f", -- $03fdc
          16349 => x"7f", -- $03fdd
          16350 => x"7f", -- $03fde
          16351 => x"7f", -- $03fdf
          16352 => x"7f", -- $03fe0
          16353 => x"7f", -- $03fe1
          16354 => x"7f", -- $03fe2
          16355 => x"7f", -- $03fe3
          16356 => x"7f", -- $03fe4
          16357 => x"7f", -- $03fe5
          16358 => x"7f", -- $03fe6
          16359 => x"7f", -- $03fe7
          16360 => x"80", -- $03fe8
          16361 => x"80", -- $03fe9
          16362 => x"80", -- $03fea
          16363 => x"80", -- $03feb
          16364 => x"80", -- $03fec
          16365 => x"80", -- $03fed
          16366 => x"80", -- $03fee
          16367 => x"80", -- $03fef
          16368 => x"80", -- $03ff0
          16369 => x"80", -- $03ff1
          16370 => x"80", -- $03ff2
          16371 => x"80", -- $03ff3
          16372 => x"80", -- $03ff4
          16373 => x"80", -- $03ff5
          16374 => x"80", -- $03ff6
          16375 => x"80", -- $03ff7
          16376 => x"7f", -- $03ff8
          16377 => x"7f", -- $03ff9
          16378 => x"80", -- $03ffa
          16379 => x"7f", -- $03ffb
          16380 => x"7f", -- $03ffc
          16381 => x"7f", -- $03ffd
          16382 => x"7f", -- $03ffe
          16383 => x"7f", -- $03fff
          16384 => x"7f", -- $04000
          16385 => x"7f", -- $04001
          16386 => x"7f", -- $04002
          16387 => x"7f", -- $04003
          16388 => x"7f", -- $04004
          16389 => x"7f", -- $04005
          16390 => x"7f", -- $04006
          16391 => x"7f", -- $04007
          16392 => x"7f", -- $04008
          16393 => x"7f", -- $04009
          16394 => x"7f", -- $0400a
          16395 => x"7f", -- $0400b
          16396 => x"7f", -- $0400c
          16397 => x"7f", -- $0400d
          16398 => x"7f", -- $0400e
          16399 => x"7f", -- $0400f
          16400 => x"7f", -- $04010
          16401 => x"7f", -- $04011
          16402 => x"7f", -- $04012
          16403 => x"7f", -- $04013
          16404 => x"7f", -- $04014
          16405 => x"7f", -- $04015
          16406 => x"7f", -- $04016
          16407 => x"7f", -- $04017
          16408 => x"7f", -- $04018
          16409 => x"7f", -- $04019
          16410 => x"7f", -- $0401a
          16411 => x"7f", -- $0401b
          16412 => x"7f", -- $0401c
          16413 => x"7f", -- $0401d
          16414 => x"7f", -- $0401e
          16415 => x"7f", -- $0401f
          16416 => x"7f", -- $04020
          16417 => x"7f", -- $04021
          16418 => x"7f", -- $04022
          16419 => x"7f", -- $04023
          16420 => x"7f", -- $04024
          16421 => x"7f", -- $04025
          16422 => x"7f", -- $04026
          16423 => x"7f", -- $04027
          16424 => x"7f", -- $04028
          16425 => x"7f", -- $04029
          16426 => x"7f", -- $0402a
          16427 => x"7f", -- $0402b
          16428 => x"7f", -- $0402c
          16429 => x"7f", -- $0402d
          16430 => x"7f", -- $0402e
          16431 => x"80", -- $0402f
          16432 => x"80", -- $04030
          16433 => x"80", -- $04031
          16434 => x"80", -- $04032
          16435 => x"80", -- $04033
          16436 => x"80", -- $04034
          16437 => x"80", -- $04035
          16438 => x"80", -- $04036
          16439 => x"80", -- $04037
          16440 => x"80", -- $04038
          16441 => x"80", -- $04039
          16442 => x"80", -- $0403a
          16443 => x"80", -- $0403b
          16444 => x"80", -- $0403c
          16445 => x"80", -- $0403d
          16446 => x"80", -- $0403e
          16447 => x"80", -- $0403f
          16448 => x"80", -- $04040
          16449 => x"80", -- $04041
          16450 => x"80", -- $04042
          16451 => x"80", -- $04043
          16452 => x"80", -- $04044
          16453 => x"80", -- $04045
          16454 => x"80", -- $04046
          16455 => x"80", -- $04047
          16456 => x"7f", -- $04048
          16457 => x"7f", -- $04049
          16458 => x"7f", -- $0404a
          16459 => x"7f", -- $0404b
          16460 => x"80", -- $0404c
          16461 => x"80", -- $0404d
          16462 => x"80", -- $0404e
          16463 => x"80", -- $0404f
          16464 => x"80", -- $04050
          16465 => x"80", -- $04051
          16466 => x"80", -- $04052
          16467 => x"80", -- $04053
          16468 => x"80", -- $04054
          16469 => x"80", -- $04055
          16470 => x"80", -- $04056
          16471 => x"80", -- $04057
          16472 => x"80", -- $04058
          16473 => x"80", -- $04059
          16474 => x"80", -- $0405a
          16475 => x"80", -- $0405b
          16476 => x"80", -- $0405c
          16477 => x"80", -- $0405d
          16478 => x"80", -- $0405e
          16479 => x"80", -- $0405f
          16480 => x"80", -- $04060
          16481 => x"80", -- $04061
          16482 => x"80", -- $04062
          16483 => x"80", -- $04063
          16484 => x"80", -- $04064
          16485 => x"80", -- $04065
          16486 => x"80", -- $04066
          16487 => x"80", -- $04067
          16488 => x"80", -- $04068
          16489 => x"80", -- $04069
          16490 => x"80", -- $0406a
          16491 => x"80", -- $0406b
          16492 => x"80", -- $0406c
          16493 => x"80", -- $0406d
          16494 => x"80", -- $0406e
          16495 => x"80", -- $0406f
          16496 => x"80", -- $04070
          16497 => x"80", -- $04071
          16498 => x"80", -- $04072
          16499 => x"80", -- $04073
          16500 => x"80", -- $04074
          16501 => x"7f", -- $04075
          16502 => x"7f", -- $04076
          16503 => x"7f", -- $04077
          16504 => x"7f", -- $04078
          16505 => x"7f", -- $04079
          16506 => x"7f", -- $0407a
          16507 => x"7f", -- $0407b
          16508 => x"7f", -- $0407c
          16509 => x"7f", -- $0407d
          16510 => x"7f", -- $0407e
          16511 => x"7f", -- $0407f
          16512 => x"7f", -- $04080
          16513 => x"7f", -- $04081
          16514 => x"7f", -- $04082
          16515 => x"7f", -- $04083
          16516 => x"7f", -- $04084
          16517 => x"7f", -- $04085
          16518 => x"7f", -- $04086
          16519 => x"7f", -- $04087
          16520 => x"7f", -- $04088
          16521 => x"7f", -- $04089
          16522 => x"7e", -- $0408a
          16523 => x"7e", -- $0408b
          16524 => x"7f", -- $0408c
          16525 => x"7f", -- $0408d
          16526 => x"7f", -- $0408e
          16527 => x"7f", -- $0408f
          16528 => x"7f", -- $04090
          16529 => x"7f", -- $04091
          16530 => x"7e", -- $04092
          16531 => x"7e", -- $04093
          16532 => x"7e", -- $04094
          16533 => x"7e", -- $04095
          16534 => x"7e", -- $04096
          16535 => x"7e", -- $04097
          16536 => x"7e", -- $04098
          16537 => x"7f", -- $04099
          16538 => x"7f", -- $0409a
          16539 => x"7e", -- $0409b
          16540 => x"7e", -- $0409c
          16541 => x"7f", -- $0409d
          16542 => x"7e", -- $0409e
          16543 => x"7e", -- $0409f
          16544 => x"7e", -- $040a0
          16545 => x"7e", -- $040a1
          16546 => x"7e", -- $040a2
          16547 => x"7c", -- $040a3
          16548 => x"7d", -- $040a4
          16549 => x"7d", -- $040a5
          16550 => x"7e", -- $040a6
          16551 => x"7d", -- $040a7
          16552 => x"7c", -- $040a8
          16553 => x"7c", -- $040a9
          16554 => x"7c", -- $040aa
          16555 => x"7c", -- $040ab
          16556 => x"7d", -- $040ac
          16557 => x"7d", -- $040ad
          16558 => x"7d", -- $040ae
          16559 => x"7d", -- $040af
          16560 => x"7e", -- $040b0
          16561 => x"7e", -- $040b1
          16562 => x"7e", -- $040b2
          16563 => x"7e", -- $040b3
          16564 => x"7f", -- $040b4
          16565 => x"7f", -- $040b5
          16566 => x"7f", -- $040b6
          16567 => x"7f", -- $040b7
          16568 => x"7f", -- $040b8
          16569 => x"7e", -- $040b9
          16570 => x"7e", -- $040ba
          16571 => x"7e", -- $040bb
          16572 => x"7e", -- $040bc
          16573 => x"7e", -- $040bd
          16574 => x"7e", -- $040be
          16575 => x"7d", -- $040bf
          16576 => x"7d", -- $040c0
          16577 => x"7e", -- $040c1
          16578 => x"7e", -- $040c2
          16579 => x"7f", -- $040c3
          16580 => x"7f", -- $040c4
          16581 => x"7e", -- $040c5
          16582 => x"7e", -- $040c6
          16583 => x"7e", -- $040c7
          16584 => x"7e", -- $040c8
          16585 => x"7f", -- $040c9
          16586 => x"7f", -- $040ca
          16587 => x"7f", -- $040cb
          16588 => x"7f", -- $040cc
          16589 => x"80", -- $040cd
          16590 => x"80", -- $040ce
          16591 => x"80", -- $040cf
          16592 => x"80", -- $040d0
          16593 => x"80", -- $040d1
          16594 => x"80", -- $040d2
          16595 => x"80", -- $040d3
          16596 => x"80", -- $040d4
          16597 => x"80", -- $040d5
          16598 => x"7f", -- $040d6
          16599 => x"7f", -- $040d7
          16600 => x"80", -- $040d8
          16601 => x"80", -- $040d9
          16602 => x"80", -- $040da
          16603 => x"80", -- $040db
          16604 => x"7f", -- $040dc
          16605 => x"7f", -- $040dd
          16606 => x"80", -- $040de
          16607 => x"80", -- $040df
          16608 => x"80", -- $040e0
          16609 => x"80", -- $040e1
          16610 => x"80", -- $040e2
          16611 => x"80", -- $040e3
          16612 => x"80", -- $040e4
          16613 => x"80", -- $040e5
          16614 => x"80", -- $040e6
          16615 => x"80", -- $040e7
          16616 => x"80", -- $040e8
          16617 => x"80", -- $040e9
          16618 => x"80", -- $040ea
          16619 => x"80", -- $040eb
          16620 => x"80", -- $040ec
          16621 => x"80", -- $040ed
          16622 => x"80", -- $040ee
          16623 => x"80", -- $040ef
          16624 => x"80", -- $040f0
          16625 => x"80", -- $040f1
          16626 => x"80", -- $040f2
          16627 => x"80", -- $040f3
          16628 => x"80", -- $040f4
          16629 => x"80", -- $040f5
          16630 => x"80", -- $040f6
          16631 => x"80", -- $040f7
          16632 => x"80", -- $040f8
          16633 => x"80", -- $040f9
          16634 => x"81", -- $040fa
          16635 => x"81", -- $040fb
          16636 => x"81", -- $040fc
          16637 => x"80", -- $040fd
          16638 => x"80", -- $040fe
          16639 => x"7f", -- $040ff
          16640 => x"80", -- $04100
          16641 => x"80", -- $04101
          16642 => x"80", -- $04102
          16643 => x"80", -- $04103
          16644 => x"80", -- $04104
          16645 => x"80", -- $04105
          16646 => x"80", -- $04106
          16647 => x"80", -- $04107
          16648 => x"80", -- $04108
          16649 => x"81", -- $04109
          16650 => x"80", -- $0410a
          16651 => x"81", -- $0410b
          16652 => x"80", -- $0410c
          16653 => x"80", -- $0410d
          16654 => x"80", -- $0410e
          16655 => x"80", -- $0410f
          16656 => x"80", -- $04110
          16657 => x"81", -- $04111
          16658 => x"81", -- $04112
          16659 => x"82", -- $04113
          16660 => x"82", -- $04114
          16661 => x"81", -- $04115
          16662 => x"80", -- $04116
          16663 => x"80", -- $04117
          16664 => x"80", -- $04118
          16665 => x"80", -- $04119
          16666 => x"80", -- $0411a
          16667 => x"80", -- $0411b
          16668 => x"80", -- $0411c
          16669 => x"80", -- $0411d
          16670 => x"80", -- $0411e
          16671 => x"80", -- $0411f
          16672 => x"80", -- $04120
          16673 => x"80", -- $04121
          16674 => x"80", -- $04122
          16675 => x"81", -- $04123
          16676 => x"82", -- $04124
          16677 => x"82", -- $04125
          16678 => x"81", -- $04126
          16679 => x"81", -- $04127
          16680 => x"81", -- $04128
          16681 => x"81", -- $04129
          16682 => x"80", -- $0412a
          16683 => x"80", -- $0412b
          16684 => x"81", -- $0412c
          16685 => x"80", -- $0412d
          16686 => x"80", -- $0412e
          16687 => x"80", -- $0412f
          16688 => x"80", -- $04130
          16689 => x"7f", -- $04131
          16690 => x"7f", -- $04132
          16691 => x"7f", -- $04133
          16692 => x"80", -- $04134
          16693 => x"80", -- $04135
          16694 => x"80", -- $04136
          16695 => x"81", -- $04137
          16696 => x"81", -- $04138
          16697 => x"81", -- $04139
          16698 => x"81", -- $0413a
          16699 => x"82", -- $0413b
          16700 => x"81", -- $0413c
          16701 => x"80", -- $0413d
          16702 => x"80", -- $0413e
          16703 => x"80", -- $0413f
          16704 => x"80", -- $04140
          16705 => x"7f", -- $04141
          16706 => x"80", -- $04142
          16707 => x"80", -- $04143
          16708 => x"80", -- $04144
          16709 => x"80", -- $04145
          16710 => x"81", -- $04146
          16711 => x"81", -- $04147
          16712 => x"81", -- $04148
          16713 => x"80", -- $04149
          16714 => x"80", -- $0414a
          16715 => x"80", -- $0414b
          16716 => x"80", -- $0414c
          16717 => x"80", -- $0414d
          16718 => x"80", -- $0414e
          16719 => x"80", -- $0414f
          16720 => x"81", -- $04150
          16721 => x"81", -- $04151
          16722 => x"81", -- $04152
          16723 => x"80", -- $04153
          16724 => x"80", -- $04154
          16725 => x"80", -- $04155
          16726 => x"80", -- $04156
          16727 => x"80", -- $04157
          16728 => x"80", -- $04158
          16729 => x"81", -- $04159
          16730 => x"81", -- $0415a
          16731 => x"82", -- $0415b
          16732 => x"81", -- $0415c
          16733 => x"81", -- $0415d
          16734 => x"80", -- $0415e
          16735 => x"80", -- $0415f
          16736 => x"80", -- $04160
          16737 => x"80", -- $04161
          16738 => x"80", -- $04162
          16739 => x"80", -- $04163
          16740 => x"80", -- $04164
          16741 => x"80", -- $04165
          16742 => x"80", -- $04166
          16743 => x"80", -- $04167
          16744 => x"80", -- $04168
          16745 => x"80", -- $04169
          16746 => x"80", -- $0416a
          16747 => x"81", -- $0416b
          16748 => x"81", -- $0416c
          16749 => x"81", -- $0416d
          16750 => x"81", -- $0416e
          16751 => x"80", -- $0416f
          16752 => x"80", -- $04170
          16753 => x"80", -- $04171
          16754 => x"80", -- $04172
          16755 => x"80", -- $04173
          16756 => x"80", -- $04174
          16757 => x"80", -- $04175
          16758 => x"80", -- $04176
          16759 => x"81", -- $04177
          16760 => x"81", -- $04178
          16761 => x"80", -- $04179
          16762 => x"80", -- $0417a
          16763 => x"80", -- $0417b
          16764 => x"81", -- $0417c
          16765 => x"80", -- $0417d
          16766 => x"80", -- $0417e
          16767 => x"81", -- $0417f
          16768 => x"80", -- $04180
          16769 => x"80", -- $04181
          16770 => x"7f", -- $04182
          16771 => x"7f", -- $04183
          16772 => x"80", -- $04184
          16773 => x"81", -- $04185
          16774 => x"82", -- $04186
          16775 => x"82", -- $04187
          16776 => x"81", -- $04188
          16777 => x"80", -- $04189
          16778 => x"80", -- $0418a
          16779 => x"80", -- $0418b
          16780 => x"80", -- $0418c
          16781 => x"80", -- $0418d
          16782 => x"81", -- $0418e
          16783 => x"82", -- $0418f
          16784 => x"82", -- $04190
          16785 => x"81", -- $04191
          16786 => x"81", -- $04192
          16787 => x"80", -- $04193
          16788 => x"80", -- $04194
          16789 => x"80", -- $04195
          16790 => x"80", -- $04196
          16791 => x"80", -- $04197
          16792 => x"80", -- $04198
          16793 => x"80", -- $04199
          16794 => x"81", -- $0419a
          16795 => x"81", -- $0419b
          16796 => x"81", -- $0419c
          16797 => x"80", -- $0419d
          16798 => x"80", -- $0419e
          16799 => x"80", -- $0419f
          16800 => x"81", -- $041a0
          16801 => x"81", -- $041a1
          16802 => x"81", -- $041a2
          16803 => x"81", -- $041a3
          16804 => x"80", -- $041a4
          16805 => x"80", -- $041a5
          16806 => x"80", -- $041a6
          16807 => x"80", -- $041a7
          16808 => x"80", -- $041a8
          16809 => x"81", -- $041a9
          16810 => x"81", -- $041aa
          16811 => x"81", -- $041ab
          16812 => x"80", -- $041ac
          16813 => x"80", -- $041ad
          16814 => x"80", -- $041ae
          16815 => x"80", -- $041af
          16816 => x"80", -- $041b0
          16817 => x"81", -- $041b1
          16818 => x"82", -- $041b2
          16819 => x"81", -- $041b3
          16820 => x"80", -- $041b4
          16821 => x"80", -- $041b5
          16822 => x"80", -- $041b6
          16823 => x"80", -- $041b7
          16824 => x"80", -- $041b8
          16825 => x"81", -- $041b9
          16826 => x"81", -- $041ba
          16827 => x"80", -- $041bb
          16828 => x"80", -- $041bc
          16829 => x"80", -- $041bd
          16830 => x"80", -- $041be
          16831 => x"81", -- $041bf
          16832 => x"81", -- $041c0
          16833 => x"82", -- $041c1
          16834 => x"82", -- $041c2
          16835 => x"81", -- $041c3
          16836 => x"80", -- $041c4
          16837 => x"80", -- $041c5
          16838 => x"80", -- $041c6
          16839 => x"80", -- $041c7
          16840 => x"81", -- $041c8
          16841 => x"81", -- $041c9
          16842 => x"81", -- $041ca
          16843 => x"81", -- $041cb
          16844 => x"80", -- $041cc
          16845 => x"80", -- $041cd
          16846 => x"81", -- $041ce
          16847 => x"81", -- $041cf
          16848 => x"81", -- $041d0
          16849 => x"81", -- $041d1
          16850 => x"81", -- $041d2
          16851 => x"80", -- $041d3
          16852 => x"80", -- $041d4
          16853 => x"80", -- $041d5
          16854 => x"80", -- $041d6
          16855 => x"81", -- $041d7
          16856 => x"81", -- $041d8
          16857 => x"81", -- $041d9
          16858 => x"80", -- $041da
          16859 => x"80", -- $041db
          16860 => x"80", -- $041dc
          16861 => x"80", -- $041dd
          16862 => x"81", -- $041de
          16863 => x"82", -- $041df
          16864 => x"82", -- $041e0
          16865 => x"82", -- $041e1
          16866 => x"82", -- $041e2
          16867 => x"81", -- $041e3
          16868 => x"80", -- $041e4
          16869 => x"7f", -- $041e5
          16870 => x"7f", -- $041e6
          16871 => x"80", -- $041e7
          16872 => x"81", -- $041e8
          16873 => x"82", -- $041e9
          16874 => x"82", -- $041ea
          16875 => x"81", -- $041eb
          16876 => x"80", -- $041ec
          16877 => x"80", -- $041ed
          16878 => x"80", -- $041ee
          16879 => x"81", -- $041ef
          16880 => x"82", -- $041f0
          16881 => x"82", -- $041f1
          16882 => x"81", -- $041f2
          16883 => x"81", -- $041f3
          16884 => x"80", -- $041f4
          16885 => x"80", -- $041f5
          16886 => x"80", -- $041f6
          16887 => x"81", -- $041f7
          16888 => x"81", -- $041f8
          16889 => x"81", -- $041f9
          16890 => x"81", -- $041fa
          16891 => x"80", -- $041fb
          16892 => x"80", -- $041fc
          16893 => x"80", -- $041fd
          16894 => x"81", -- $041fe
          16895 => x"82", -- $041ff
          16896 => x"81", -- $04200
          16897 => x"81", -- $04201
          16898 => x"80", -- $04202
          16899 => x"7f", -- $04203
          16900 => x"7f", -- $04204
          16901 => x"80", -- $04205
          16902 => x"81", -- $04206
          16903 => x"82", -- $04207
          16904 => x"82", -- $04208
          16905 => x"81", -- $04209
          16906 => x"80", -- $0420a
          16907 => x"80", -- $0420b
          16908 => x"80", -- $0420c
          16909 => x"81", -- $0420d
          16910 => x"81", -- $0420e
          16911 => x"82", -- $0420f
          16912 => x"82", -- $04210
          16913 => x"81", -- $04211
          16914 => x"81", -- $04212
          16915 => x"80", -- $04213
          16916 => x"80", -- $04214
          16917 => x"80", -- $04215
          16918 => x"80", -- $04216
          16919 => x"80", -- $04217
          16920 => x"80", -- $04218
          16921 => x"80", -- $04219
          16922 => x"80", -- $0421a
          16923 => x"80", -- $0421b
          16924 => x"81", -- $0421c
          16925 => x"81", -- $0421d
          16926 => x"82", -- $0421e
          16927 => x"81", -- $0421f
          16928 => x"81", -- $04220
          16929 => x"81", -- $04221
          16930 => x"81", -- $04222
          16931 => x"81", -- $04223
          16932 => x"82", -- $04224
          16933 => x"82", -- $04225
          16934 => x"81", -- $04226
          16935 => x"80", -- $04227
          16936 => x"80", -- $04228
          16937 => x"80", -- $04229
          16938 => x"80", -- $0422a
          16939 => x"80", -- $0422b
          16940 => x"81", -- $0422c
          16941 => x"81", -- $0422d
          16942 => x"81", -- $0422e
          16943 => x"81", -- $0422f
          16944 => x"81", -- $04230
          16945 => x"81", -- $04231
          16946 => x"81", -- $04232
          16947 => x"81", -- $04233
          16948 => x"80", -- $04234
          16949 => x"80", -- $04235
          16950 => x"80", -- $04236
          16951 => x"80", -- $04237
          16952 => x"81", -- $04238
          16953 => x"81", -- $04239
          16954 => x"80", -- $0423a
          16955 => x"80", -- $0423b
          16956 => x"80", -- $0423c
          16957 => x"80", -- $0423d
          16958 => x"80", -- $0423e
          16959 => x"80", -- $0423f
          16960 => x"81", -- $04240
          16961 => x"81", -- $04241
          16962 => x"81", -- $04242
          16963 => x"80", -- $04243
          16964 => x"80", -- $04244
          16965 => x"80", -- $04245
          16966 => x"80", -- $04246
          16967 => x"81", -- $04247
          16968 => x"81", -- $04248
          16969 => x"81", -- $04249
          16970 => x"80", -- $0424a
          16971 => x"80", -- $0424b
          16972 => x"80", -- $0424c
          16973 => x"80", -- $0424d
          16974 => x"80", -- $0424e
          16975 => x"81", -- $0424f
          16976 => x"80", -- $04250
          16977 => x"80", -- $04251
          16978 => x"80", -- $04252
          16979 => x"80", -- $04253
          16980 => x"80", -- $04254
          16981 => x"80", -- $04255
          16982 => x"80", -- $04256
          16983 => x"80", -- $04257
          16984 => x"80", -- $04258
          16985 => x"80", -- $04259
          16986 => x"80", -- $0425a
          16987 => x"80", -- $0425b
          16988 => x"80", -- $0425c
          16989 => x"80", -- $0425d
          16990 => x"80", -- $0425e
          16991 => x"80", -- $0425f
          16992 => x"80", -- $04260
          16993 => x"80", -- $04261
          16994 => x"80", -- $04262
          16995 => x"80", -- $04263
          16996 => x"80", -- $04264
          16997 => x"7f", -- $04265
          16998 => x"7f", -- $04266
          16999 => x"7f", -- $04267
          17000 => x"7e", -- $04268
          17001 => x"7e", -- $04269
          17002 => x"7f", -- $0426a
          17003 => x"7f", -- $0426b
          17004 => x"80", -- $0426c
          17005 => x"7f", -- $0426d
          17006 => x"7e", -- $0426e
          17007 => x"7e", -- $0426f
          17008 => x"7e", -- $04270
          17009 => x"7f", -- $04271
          17010 => x"7f", -- $04272
          17011 => x"7f", -- $04273
          17012 => x"7f", -- $04274
          17013 => x"7f", -- $04275
          17014 => x"7e", -- $04276
          17015 => x"7e", -- $04277
          17016 => x"7e", -- $04278
          17017 => x"7f", -- $04279
          17018 => x"7f", -- $0427a
          17019 => x"80", -- $0427b
          17020 => x"80", -- $0427c
          17021 => x"7f", -- $0427d
          17022 => x"7f", -- $0427e
          17023 => x"80", -- $0427f
          17024 => x"80", -- $04280
          17025 => x"81", -- $04281
          17026 => x"82", -- $04282
          17027 => x"82", -- $04283
          17028 => x"82", -- $04284
          17029 => x"83", -- $04285
          17030 => x"84", -- $04286
          17031 => x"84", -- $04287
          17032 => x"84", -- $04288
          17033 => x"84", -- $04289
          17034 => x"84", -- $0428a
          17035 => x"85", -- $0428b
          17036 => x"86", -- $0428c
          17037 => x"86", -- $0428d
          17038 => x"86", -- $0428e
          17039 => x"85", -- $0428f
          17040 => x"86", -- $04290
          17041 => x"86", -- $04291
          17042 => x"87", -- $04292
          17043 => x"87", -- $04293
          17044 => x"87", -- $04294
          17045 => x"87", -- $04295
          17046 => x"88", -- $04296
          17047 => x"88", -- $04297
          17048 => x"87", -- $04298
          17049 => x"87", -- $04299
          17050 => x"87", -- $0429a
          17051 => x"86", -- $0429b
          17052 => x"85", -- $0429c
          17053 => x"85", -- $0429d
          17054 => x"84", -- $0429e
          17055 => x"83", -- $0429f
          17056 => x"82", -- $042a0
          17057 => x"82", -- $042a1
          17058 => x"81", -- $042a2
          17059 => x"81", -- $042a3
          17060 => x"80", -- $042a4
          17061 => x"80", -- $042a5
          17062 => x"80", -- $042a6
          17063 => x"80", -- $042a7
          17064 => x"80", -- $042a8
          17065 => x"7f", -- $042a9
          17066 => x"7f", -- $042aa
          17067 => x"7e", -- $042ab
          17068 => x"7e", -- $042ac
          17069 => x"7d", -- $042ad
          17070 => x"7c", -- $042ae
          17071 => x"7b", -- $042af
          17072 => x"7a", -- $042b0
          17073 => x"7a", -- $042b1
          17074 => x"79", -- $042b2
          17075 => x"79", -- $042b3
          17076 => x"79", -- $042b4
          17077 => x"79", -- $042b5
          17078 => x"78", -- $042b6
          17079 => x"78", -- $042b7
          17080 => x"78", -- $042b8
          17081 => x"78", -- $042b9
          17082 => x"78", -- $042ba
          17083 => x"78", -- $042bb
          17084 => x"78", -- $042bc
          17085 => x"78", -- $042bd
          17086 => x"78", -- $042be
          17087 => x"77", -- $042bf
          17088 => x"77", -- $042c0
          17089 => x"77", -- $042c1
          17090 => x"77", -- $042c2
          17091 => x"77", -- $042c3
          17092 => x"78", -- $042c4
          17093 => x"77", -- $042c5
          17094 => x"76", -- $042c6
          17095 => x"76", -- $042c7
          17096 => x"76", -- $042c8
          17097 => x"77", -- $042c9
          17098 => x"78", -- $042ca
          17099 => x"79", -- $042cb
          17100 => x"79", -- $042cc
          17101 => x"78", -- $042cd
          17102 => x"78", -- $042ce
          17103 => x"79", -- $042cf
          17104 => x"7a", -- $042d0
          17105 => x"7b", -- $042d1
          17106 => x"7b", -- $042d2
          17107 => x"7b", -- $042d3
          17108 => x"7b", -- $042d4
          17109 => x"7c", -- $042d5
          17110 => x"7c", -- $042d6
          17111 => x"7d", -- $042d7
          17112 => x"7d", -- $042d8
          17113 => x"7e", -- $042d9
          17114 => x"7f", -- $042da
          17115 => x"7f", -- $042db
          17116 => x"80", -- $042dc
          17117 => x"80", -- $042dd
          17118 => x"80", -- $042de
          17119 => x"80", -- $042df
          17120 => x"81", -- $042e0
          17121 => x"83", -- $042e1
          17122 => x"84", -- $042e2
          17123 => x"85", -- $042e3
          17124 => x"85", -- $042e4
          17125 => x"85", -- $042e5
          17126 => x"86", -- $042e6
          17127 => x"86", -- $042e7
          17128 => x"87", -- $042e8
          17129 => x"88", -- $042e9
          17130 => x"88", -- $042ea
          17131 => x"88", -- $042eb
          17132 => x"89", -- $042ec
          17133 => x"89", -- $042ed
          17134 => x"8a", -- $042ee
          17135 => x"8a", -- $042ef
          17136 => x"8a", -- $042f0
          17137 => x"8a", -- $042f1
          17138 => x"8b", -- $042f2
          17139 => x"8b", -- $042f3
          17140 => x"8a", -- $042f4
          17141 => x"8a", -- $042f5
          17142 => x"8a", -- $042f6
          17143 => x"8a", -- $042f7
          17144 => x"8a", -- $042f8
          17145 => x"8a", -- $042f9
          17146 => x"89", -- $042fa
          17147 => x"89", -- $042fb
          17148 => x"88", -- $042fc
          17149 => x"88", -- $042fd
          17150 => x"88", -- $042fe
          17151 => x"87", -- $042ff
          17152 => x"87", -- $04300
          17153 => x"87", -- $04301
          17154 => x"86", -- $04302
          17155 => x"85", -- $04303
          17156 => x"85", -- $04304
          17157 => x"84", -- $04305
          17158 => x"83", -- $04306
          17159 => x"83", -- $04307
          17160 => x"82", -- $04308
          17161 => x"82", -- $04309
          17162 => x"81", -- $0430a
          17163 => x"80", -- $0430b
          17164 => x"80", -- $0430c
          17165 => x"80", -- $0430d
          17166 => x"80", -- $0430e
          17167 => x"7f", -- $0430f
          17168 => x"7e", -- $04310
          17169 => x"7e", -- $04311
          17170 => x"7e", -- $04312
          17171 => x"7e", -- $04313
          17172 => x"7e", -- $04314
          17173 => x"7d", -- $04315
          17174 => x"7c", -- $04316
          17175 => x"7c", -- $04317
          17176 => x"7c", -- $04318
          17177 => x"7d", -- $04319
          17178 => x"7c", -- $0431a
          17179 => x"7c", -- $0431b
          17180 => x"7b", -- $0431c
          17181 => x"7b", -- $0431d
          17182 => x"7b", -- $0431e
          17183 => x"7b", -- $0431f
          17184 => x"7b", -- $04320
          17185 => x"7b", -- $04321
          17186 => x"7b", -- $04322
          17187 => x"7b", -- $04323
          17188 => x"7b", -- $04324
          17189 => x"7a", -- $04325
          17190 => x"7a", -- $04326
          17191 => x"7a", -- $04327
          17192 => x"7a", -- $04328
          17193 => x"7a", -- $04329
          17194 => x"7a", -- $0432a
          17195 => x"7a", -- $0432b
          17196 => x"79", -- $0432c
          17197 => x"78", -- $0432d
          17198 => x"78", -- $0432e
          17199 => x"77", -- $0432f
          17200 => x"78", -- $04330
          17201 => x"78", -- $04331
          17202 => x"78", -- $04332
          17203 => x"78", -- $04333
          17204 => x"78", -- $04334
          17205 => x"78", -- $04335
          17206 => x"78", -- $04336
          17207 => x"79", -- $04337
          17208 => x"7a", -- $04338
          17209 => x"7a", -- $04339
          17210 => x"7a", -- $0433a
          17211 => x"7b", -- $0433b
          17212 => x"7b", -- $0433c
          17213 => x"7c", -- $0433d
          17214 => x"7c", -- $0433e
          17215 => x"7d", -- $0433f
          17216 => x"7f", -- $04340
          17217 => x"80", -- $04341
          17218 => x"80", -- $04342
          17219 => x"81", -- $04343
          17220 => x"81", -- $04344
          17221 => x"81", -- $04345
          17222 => x"82", -- $04346
          17223 => x"84", -- $04347
          17224 => x"86", -- $04348
          17225 => x"86", -- $04349
          17226 => x"86", -- $0434a
          17227 => x"86", -- $0434b
          17228 => x"85", -- $0434c
          17229 => x"86", -- $0434d
          17230 => x"86", -- $0434e
          17231 => x"86", -- $0434f
          17232 => x"85", -- $04350
          17233 => x"85", -- $04351
          17234 => x"84", -- $04352
          17235 => x"83", -- $04353
          17236 => x"82", -- $04354
          17237 => x"82", -- $04355
          17238 => x"83", -- $04356
          17239 => x"83", -- $04357
          17240 => x"82", -- $04358
          17241 => x"80", -- $04359
          17242 => x"7f", -- $0435a
          17243 => x"7d", -- $0435b
          17244 => x"7c", -- $0435c
          17245 => x"7d", -- $0435d
          17246 => x"7e", -- $0435e
          17247 => x"7f", -- $0435f
          17248 => x"80", -- $04360
          17249 => x"80", -- $04361
          17250 => x"82", -- $04362
          17251 => x"83", -- $04363
          17252 => x"85", -- $04364
          17253 => x"87", -- $04365
          17254 => x"89", -- $04366
          17255 => x"88", -- $04367
          17256 => x"87", -- $04368
          17257 => x"86", -- $04369
          17258 => x"87", -- $0436a
          17259 => x"89", -- $0436b
          17260 => x"8c", -- $0436c
          17261 => x"8d", -- $0436d
          17262 => x"8d", -- $0436e
          17263 => x"8c", -- $0436f
          17264 => x"8b", -- $04370
          17265 => x"88", -- $04371
          17266 => x"85", -- $04372
          17267 => x"83", -- $04373
          17268 => x"83", -- $04374
          17269 => x"85", -- $04375
          17270 => x"86", -- $04376
          17271 => x"85", -- $04377
          17272 => x"81", -- $04378
          17273 => x"7f", -- $04379
          17274 => x"7e", -- $0437a
          17275 => x"7e", -- $0437b
          17276 => x"7d", -- $0437c
          17277 => x"7a", -- $0437d
          17278 => x"76", -- $0437e
          17279 => x"73", -- $0437f
          17280 => x"72", -- $04380
          17281 => x"71", -- $04381
          17282 => x"72", -- $04382
          17283 => x"73", -- $04383
          17284 => x"77", -- $04384
          17285 => x"7b", -- $04385
          17286 => x"7e", -- $04386
          17287 => x"7f", -- $04387
          17288 => x"7d", -- $04388
          17289 => x"7d", -- $04389
          17290 => x"7d", -- $0438a
          17291 => x"7d", -- $0438b
          17292 => x"7c", -- $0438c
          17293 => x"7c", -- $0438d
          17294 => x"7c", -- $0438e
          17295 => x"7d", -- $0438f
          17296 => x"7f", -- $04390
          17297 => x"80", -- $04391
          17298 => x"80", -- $04392
          17299 => x"81", -- $04393
          17300 => x"82", -- $04394
          17301 => x"83", -- $04395
          17302 => x"83", -- $04396
          17303 => x"81", -- $04397
          17304 => x"80", -- $04398
          17305 => x"7f", -- $04399
          17306 => x"7e", -- $0439a
          17307 => x"7e", -- $0439b
          17308 => x"7e", -- $0439c
          17309 => x"7e", -- $0439d
          17310 => x"7e", -- $0439e
          17311 => x"7f", -- $0439f
          17312 => x"7f", -- $043a0
          17313 => x"7e", -- $043a1
          17314 => x"7b", -- $043a2
          17315 => x"76", -- $043a3
          17316 => x"72", -- $043a4
          17317 => x"6e", -- $043a5
          17318 => x"6c", -- $043a6
          17319 => x"6d", -- $043a7
          17320 => x"6f", -- $043a8
          17321 => x"74", -- $043a9
          17322 => x"78", -- $043aa
          17323 => x"7c", -- $043ab
          17324 => x"7e", -- $043ac
          17325 => x"7f", -- $043ad
          17326 => x"7f", -- $043ae
          17327 => x"7f", -- $043af
          17328 => x"7e", -- $043b0
          17329 => x"7e", -- $043b1
          17330 => x"7e", -- $043b2
          17331 => x"7f", -- $043b3
          17332 => x"7f", -- $043b4
          17333 => x"80", -- $043b5
          17334 => x"81", -- $043b6
          17335 => x"82", -- $043b7
          17336 => x"84", -- $043b8
          17337 => x"84", -- $043b9
          17338 => x"84", -- $043ba
          17339 => x"83", -- $043bb
          17340 => x"84", -- $043bc
          17341 => x"85", -- $043bd
          17342 => x"86", -- $043be
          17343 => x"88", -- $043bf
          17344 => x"89", -- $043c0
          17345 => x"89", -- $043c1
          17346 => x"89", -- $043c2
          17347 => x"88", -- $043c3
          17348 => x"87", -- $043c4
          17349 => x"86", -- $043c5
          17350 => x"84", -- $043c6
          17351 => x"82", -- $043c7
          17352 => x"80", -- $043c8
          17353 => x"7d", -- $043c9
          17354 => x"7b", -- $043ca
          17355 => x"7b", -- $043cb
          17356 => x"7d", -- $043cc
          17357 => x"7f", -- $043cd
          17358 => x"80", -- $043ce
          17359 => x"81", -- $043cf
          17360 => x"80", -- $043d0
          17361 => x"7e", -- $043d1
          17362 => x"7a", -- $043d2
          17363 => x"77", -- $043d3
          17364 => x"76", -- $043d4
          17365 => x"76", -- $043d5
          17366 => x"78", -- $043d6
          17367 => x"7b", -- $043d7
          17368 => x"7d", -- $043d8
          17369 => x"80", -- $043d9
          17370 => x"81", -- $043da
          17371 => x"83", -- $043db
          17372 => x"84", -- $043dc
          17373 => x"84", -- $043dd
          17374 => x"85", -- $043de
          17375 => x"86", -- $043df
          17376 => x"87", -- $043e0
          17377 => x"88", -- $043e1
          17378 => x"88", -- $043e2
          17379 => x"89", -- $043e3
          17380 => x"89", -- $043e4
          17381 => x"89", -- $043e5
          17382 => x"87", -- $043e6
          17383 => x"86", -- $043e7
          17384 => x"85", -- $043e8
          17385 => x"83", -- $043e9
          17386 => x"81", -- $043ea
          17387 => x"80", -- $043eb
          17388 => x"80", -- $043ec
          17389 => x"81", -- $043ed
          17390 => x"81", -- $043ee
          17391 => x"82", -- $043ef
          17392 => x"83", -- $043f0
          17393 => x"84", -- $043f1
          17394 => x"83", -- $043f2
          17395 => x"80", -- $043f3
          17396 => x"7c", -- $043f4
          17397 => x"78", -- $043f5
          17398 => x"73", -- $043f6
          17399 => x"6f", -- $043f7
          17400 => x"6b", -- $043f8
          17401 => x"6b", -- $043f9
          17402 => x"6e", -- $043fa
          17403 => x"72", -- $043fb
          17404 => x"76", -- $043fc
          17405 => x"7b", -- $043fd
          17406 => x"7f", -- $043fe
          17407 => x"81", -- $043ff
          17408 => x"82", -- $04400
          17409 => x"80", -- $04401
          17410 => x"80", -- $04402
          17411 => x"80", -- $04403
          17412 => x"80", -- $04404
          17413 => x"80", -- $04405
          17414 => x"81", -- $04406
          17415 => x"82", -- $04407
          17416 => x"84", -- $04408
          17417 => x"84", -- $04409
          17418 => x"83", -- $0440a
          17419 => x"82", -- $0440b
          17420 => x"81", -- $0440c
          17421 => x"82", -- $0440d
          17422 => x"82", -- $0440e
          17423 => x"83", -- $0440f
          17424 => x"85", -- $04410
          17425 => x"88", -- $04411
          17426 => x"89", -- $04412
          17427 => x"89", -- $04413
          17428 => x"88", -- $04414
          17429 => x"87", -- $04415
          17430 => x"85", -- $04416
          17431 => x"83", -- $04417
          17432 => x"80", -- $04418
          17433 => x"80", -- $04419
          17434 => x"7d", -- $0441a
          17435 => x"7b", -- $0441b
          17436 => x"79", -- $0441c
          17437 => x"79", -- $0441d
          17438 => x"79", -- $0441e
          17439 => x"7b", -- $0441f
          17440 => x"7d", -- $04420
          17441 => x"7f", -- $04421
          17442 => x"80", -- $04422
          17443 => x"80", -- $04423
          17444 => x"80", -- $04424
          17445 => x"7e", -- $04425
          17446 => x"7b", -- $04426
          17447 => x"7a", -- $04427
          17448 => x"79", -- $04428
          17449 => x"79", -- $04429
          17450 => x"7c", -- $0442a
          17451 => x"7e", -- $0442b
          17452 => x"81", -- $0442c
          17453 => x"83", -- $0442d
          17454 => x"86", -- $0442e
          17455 => x"88", -- $0442f
          17456 => x"88", -- $04430
          17457 => x"88", -- $04431
          17458 => x"88", -- $04432
          17459 => x"89", -- $04433
          17460 => x"89", -- $04434
          17461 => x"89", -- $04435
          17462 => x"8a", -- $04436
          17463 => x"8c", -- $04437
          17464 => x"8c", -- $04438
          17465 => x"8c", -- $04439
          17466 => x"8b", -- $0443a
          17467 => x"8a", -- $0443b
          17468 => x"88", -- $0443c
          17469 => x"85", -- $0443d
          17470 => x"81", -- $0443e
          17471 => x"80", -- $0443f
          17472 => x"80", -- $04440
          17473 => x"80", -- $04441
          17474 => x"80", -- $04442
          17475 => x"80", -- $04443
          17476 => x"82", -- $04444
          17477 => x"82", -- $04445
          17478 => x"80", -- $04446
          17479 => x"7f", -- $04447
          17480 => x"7d", -- $04448
          17481 => x"79", -- $04449
          17482 => x"74", -- $0444a
          17483 => x"70", -- $0444b
          17484 => x"6e", -- $0444c
          17485 => x"6e", -- $0444d
          17486 => x"70", -- $0444e
          17487 => x"73", -- $0444f
          17488 => x"79", -- $04450
          17489 => x"7e", -- $04451
          17490 => x"82", -- $04452
          17491 => x"84", -- $04453
          17492 => x"85", -- $04454
          17493 => x"85", -- $04455
          17494 => x"84", -- $04456
          17495 => x"83", -- $04457
          17496 => x"83", -- $04458
          17497 => x"83", -- $04459
          17498 => x"84", -- $0445a
          17499 => x"84", -- $0445b
          17500 => x"85", -- $0445c
          17501 => x"85", -- $0445d
          17502 => x"84", -- $0445e
          17503 => x"82", -- $0445f
          17504 => x"81", -- $04460
          17505 => x"81", -- $04461
          17506 => x"81", -- $04462
          17507 => x"81", -- $04463
          17508 => x"83", -- $04464
          17509 => x"85", -- $04465
          17510 => x"86", -- $04466
          17511 => x"86", -- $04467
          17512 => x"85", -- $04468
          17513 => x"83", -- $04469
          17514 => x"81", -- $0446a
          17515 => x"7f", -- $0446b
          17516 => x"7d", -- $0446c
          17517 => x"7c", -- $0446d
          17518 => x"7b", -- $0446e
          17519 => x"7a", -- $0446f
          17520 => x"79", -- $04470
          17521 => x"79", -- $04471
          17522 => x"78", -- $04472
          17523 => x"79", -- $04473
          17524 => x"7a", -- $04474
          17525 => x"7c", -- $04475
          17526 => x"7d", -- $04476
          17527 => x"7f", -- $04477
          17528 => x"80", -- $04478
          17529 => x"80", -- $04479
          17530 => x"80", -- $0447a
          17531 => x"7f", -- $0447b
          17532 => x"7d", -- $0447c
          17533 => x"7d", -- $0447d
          17534 => x"7d", -- $0447e
          17535 => x"7f", -- $0447f
          17536 => x"81", -- $04480
          17537 => x"84", -- $04481
          17538 => x"87", -- $04482
          17539 => x"89", -- $04483
          17540 => x"8a", -- $04484
          17541 => x"8a", -- $04485
          17542 => x"89", -- $04486
          17543 => x"88", -- $04487
          17544 => x"87", -- $04488
          17545 => x"87", -- $04489
          17546 => x"87", -- $0448a
          17547 => x"87", -- $0448b
          17548 => x"88", -- $0448c
          17549 => x"88", -- $0448d
          17550 => x"87", -- $0448e
          17551 => x"86", -- $0448f
          17552 => x"85", -- $04490
          17553 => x"83", -- $04491
          17554 => x"82", -- $04492
          17555 => x"81", -- $04493
          17556 => x"81", -- $04494
          17557 => x"81", -- $04495
          17558 => x"81", -- $04496
          17559 => x"81", -- $04497
          17560 => x"81", -- $04498
          17561 => x"81", -- $04499
          17562 => x"80", -- $0449a
          17563 => x"80", -- $0449b
          17564 => x"80", -- $0449c
          17565 => x"80", -- $0449d
          17566 => x"80", -- $0449e
          17567 => x"7e", -- $0449f
          17568 => x"7c", -- $044a0
          17569 => x"7a", -- $044a1
          17570 => x"77", -- $044a2
          17571 => x"77", -- $044a3
          17572 => x"77", -- $044a4
          17573 => x"7a", -- $044a5
          17574 => x"7e", -- $044a6
          17575 => x"81", -- $044a7
          17576 => x"86", -- $044a8
          17577 => x"89", -- $044a9
          17578 => x"8a", -- $044aa
          17579 => x"89", -- $044ab
          17580 => x"87", -- $044ac
          17581 => x"85", -- $044ad
          17582 => x"83", -- $044ae
          17583 => x"81", -- $044af
          17584 => x"80", -- $044b0
          17585 => x"80", -- $044b1
          17586 => x"80", -- $044b2
          17587 => x"81", -- $044b3
          17588 => x"81", -- $044b4
          17589 => x"80", -- $044b5
          17590 => x"80", -- $044b6
          17591 => x"7e", -- $044b7
          17592 => x"7d", -- $044b8
          17593 => x"7b", -- $044b9
          17594 => x"7b", -- $044ba
          17595 => x"7c", -- $044bb
          17596 => x"7e", -- $044bc
          17597 => x"7f", -- $044bd
          17598 => x"80", -- $044be
          17599 => x"80", -- $044bf
          17600 => x"80", -- $044c0
          17601 => x"7e", -- $044c1
          17602 => x"7d", -- $044c2
          17603 => x"7c", -- $044c3
          17604 => x"7c", -- $044c4
          17605 => x"7c", -- $044c5
          17606 => x"7c", -- $044c6
          17607 => x"7d", -- $044c7
          17608 => x"7d", -- $044c8
          17609 => x"7d", -- $044c9
          17610 => x"7e", -- $044ca
          17611 => x"7f", -- $044cb
          17612 => x"80", -- $044cc
          17613 => x"82", -- $044cd
          17614 => x"84", -- $044ce
          17615 => x"85", -- $044cf
          17616 => x"84", -- $044d0
          17617 => x"83", -- $044d1
          17618 => x"80", -- $044d2
          17619 => x"7e", -- $044d3
          17620 => x"7b", -- $044d4
          17621 => x"79", -- $044d5
          17622 => x"78", -- $044d6
          17623 => x"78", -- $044d7
          17624 => x"79", -- $044d8
          17625 => x"7b", -- $044d9
          17626 => x"7d", -- $044da
          17627 => x"7f", -- $044db
          17628 => x"80", -- $044dc
          17629 => x"80", -- $044dd
          17630 => x"80", -- $044de
          17631 => x"7e", -- $044df
          17632 => x"7d", -- $044e0
          17633 => x"7c", -- $044e1
          17634 => x"7b", -- $044e2
          17635 => x"7a", -- $044e3
          17636 => x"7a", -- $044e4
          17637 => x"7a", -- $044e5
          17638 => x"7a", -- $044e6
          17639 => x"7b", -- $044e7
          17640 => x"7b", -- $044e8
          17641 => x"7c", -- $044e9
          17642 => x"7d", -- $044ea
          17643 => x"7e", -- $044eb
          17644 => x"80", -- $044ec
          17645 => x"81", -- $044ed
          17646 => x"83", -- $044ee
          17647 => x"84", -- $044ef
          17648 => x"86", -- $044f0
          17649 => x"87", -- $044f1
          17650 => x"88", -- $044f2
          17651 => x"88", -- $044f3
          17652 => x"88", -- $044f4
          17653 => x"86", -- $044f5
          17654 => x"85", -- $044f6
          17655 => x"83", -- $044f7
          17656 => x"82", -- $044f8
          17657 => x"81", -- $044f9
          17658 => x"81", -- $044fa
          17659 => x"82", -- $044fb
          17660 => x"84", -- $044fc
          17661 => x"85", -- $044fd
          17662 => x"86", -- $044fe
          17663 => x"85", -- $044ff
          17664 => x"84", -- $04500
          17665 => x"83", -- $04501
          17666 => x"81", -- $04502
          17667 => x"7f", -- $04503
          17668 => x"7d", -- $04504
          17669 => x"7c", -- $04505
          17670 => x"7b", -- $04506
          17671 => x"7a", -- $04507
          17672 => x"7a", -- $04508
          17673 => x"7b", -- $04509
          17674 => x"7c", -- $0450a
          17675 => x"7d", -- $0450b
          17676 => x"7e", -- $0450c
          17677 => x"7f", -- $0450d
          17678 => x"7f", -- $0450e
          17679 => x"7f", -- $0450f
          17680 => x"80", -- $04510
          17681 => x"80", -- $04511
          17682 => x"80", -- $04512
          17683 => x"80", -- $04513
          17684 => x"80", -- $04514
          17685 => x"80", -- $04515
          17686 => x"80", -- $04516
          17687 => x"7f", -- $04517
          17688 => x"7f", -- $04518
          17689 => x"80", -- $04519
          17690 => x"80", -- $0451a
          17691 => x"80", -- $0451b
          17692 => x"81", -- $0451c
          17693 => x"83", -- $0451d
          17694 => x"84", -- $0451e
          17695 => x"85", -- $0451f
          17696 => x"86", -- $04520
          17697 => x"87", -- $04521
          17698 => x"87", -- $04522
          17699 => x"87", -- $04523
          17700 => x"87", -- $04524
          17701 => x"86", -- $04525
          17702 => x"86", -- $04526
          17703 => x"85", -- $04527
          17704 => x"84", -- $04528
          17705 => x"82", -- $04529
          17706 => x"80", -- $0452a
          17707 => x"80", -- $0452b
          17708 => x"7f", -- $0452c
          17709 => x"7f", -- $0452d
          17710 => x"7f", -- $0452e
          17711 => x"7f", -- $0452f
          17712 => x"80", -- $04530
          17713 => x"80", -- $04531
          17714 => x"80", -- $04532
          17715 => x"7f", -- $04533
          17716 => x"7e", -- $04534
          17717 => x"7d", -- $04535
          17718 => x"7b", -- $04536
          17719 => x"7a", -- $04537
          17720 => x"79", -- $04538
          17721 => x"79", -- $04539
          17722 => x"79", -- $0453a
          17723 => x"79", -- $0453b
          17724 => x"7a", -- $0453c
          17725 => x"7b", -- $0453d
          17726 => x"7c", -- $0453e
          17727 => x"7e", -- $0453f
          17728 => x"7f", -- $04540
          17729 => x"80", -- $04541
          17730 => x"81", -- $04542
          17731 => x"82", -- $04543
          17732 => x"82", -- $04544
          17733 => x"82", -- $04545
          17734 => x"82", -- $04546
          17735 => x"81", -- $04547
          17736 => x"81", -- $04548
          17737 => x"80", -- $04549
          17738 => x"80", -- $0454a
          17739 => x"80", -- $0454b
          17740 => x"80", -- $0454c
          17741 => x"81", -- $0454d
          17742 => x"81", -- $0454e
          17743 => x"81", -- $0454f
          17744 => x"81", -- $04550
          17745 => x"81", -- $04551
          17746 => x"82", -- $04552
          17747 => x"82", -- $04553
          17748 => x"82", -- $04554
          17749 => x"82", -- $04555
          17750 => x"82", -- $04556
          17751 => x"81", -- $04557
          17752 => x"81", -- $04558
          17753 => x"81", -- $04559
          17754 => x"81", -- $0455a
          17755 => x"81", -- $0455b
          17756 => x"81", -- $0455c
          17757 => x"81", -- $0455d
          17758 => x"81", -- $0455e
          17759 => x"81", -- $0455f
          17760 => x"82", -- $04560
          17761 => x"83", -- $04561
          17762 => x"83", -- $04562
          17763 => x"84", -- $04563
          17764 => x"84", -- $04564
          17765 => x"85", -- $04565
          17766 => x"85", -- $04566
          17767 => x"85", -- $04567
          17768 => x"84", -- $04568
          17769 => x"83", -- $04569
          17770 => x"83", -- $0456a
          17771 => x"82", -- $0456b
          17772 => x"81", -- $0456c
          17773 => x"81", -- $0456d
          17774 => x"80", -- $0456e
          17775 => x"80", -- $0456f
          17776 => x"80", -- $04570
          17777 => x"80", -- $04571
          17778 => x"80", -- $04572
          17779 => x"80", -- $04573
          17780 => x"80", -- $04574
          17781 => x"80", -- $04575
          17782 => x"80", -- $04576
          17783 => x"80", -- $04577
          17784 => x"80", -- $04578
          17785 => x"80", -- $04579
          17786 => x"7f", -- $0457a
          17787 => x"7f", -- $0457b
          17788 => x"7f", -- $0457c
          17789 => x"7f", -- $0457d
          17790 => x"7f", -- $0457e
          17791 => x"7f", -- $0457f
          17792 => x"7f", -- $04580
          17793 => x"7f", -- $04581
          17794 => x"80", -- $04582
          17795 => x"80", -- $04583
          17796 => x"80", -- $04584
          17797 => x"80", -- $04585
          17798 => x"80", -- $04586
          17799 => x"7f", -- $04587
          17800 => x"7f", -- $04588
          17801 => x"7f", -- $04589
          17802 => x"7f", -- $0458a
          17803 => x"7f", -- $0458b
          17804 => x"7f", -- $0458c
          17805 => x"7f", -- $0458d
          17806 => x"7f", -- $0458e
          17807 => x"80", -- $0458f
          17808 => x"80", -- $04590
          17809 => x"80", -- $04591
          17810 => x"81", -- $04592
          17811 => x"81", -- $04593
          17812 => x"81", -- $04594
          17813 => x"81", -- $04595
          17814 => x"81", -- $04596
          17815 => x"81", -- $04597
          17816 => x"81", -- $04598
          17817 => x"81", -- $04599
          17818 => x"80", -- $0459a
          17819 => x"80", -- $0459b
          17820 => x"80", -- $0459c
          17821 => x"7f", -- $0459d
          17822 => x"7f", -- $0459e
          17823 => x"7e", -- $0459f
          17824 => x"7d", -- $045a0
          17825 => x"7d", -- $045a1
          17826 => x"7d", -- $045a2
          17827 => x"7d", -- $045a3
          17828 => x"7d", -- $045a4
          17829 => x"7d", -- $045a5
          17830 => x"7d", -- $045a6
          17831 => x"7e", -- $045a7
          17832 => x"7e", -- $045a8
          17833 => x"7e", -- $045a9
          17834 => x"7e", -- $045aa
          17835 => x"7e", -- $045ab
          17836 => x"7e", -- $045ac
          17837 => x"7e", -- $045ad
          17838 => x"7f", -- $045ae
          17839 => x"7f", -- $045af
          17840 => x"7f", -- $045b0
          17841 => x"80", -- $045b1
          17842 => x"80", -- $045b2
          17843 => x"80", -- $045b3
          17844 => x"80", -- $045b4
          17845 => x"80", -- $045b5
          17846 => x"80", -- $045b6
          17847 => x"81", -- $045b7
          17848 => x"81", -- $045b8
          17849 => x"81", -- $045b9
          17850 => x"81", -- $045ba
          17851 => x"81", -- $045bb
          17852 => x"81", -- $045bc
          17853 => x"81", -- $045bd
          17854 => x"80", -- $045be
          17855 => x"80", -- $045bf
          17856 => x"80", -- $045c0
          17857 => x"80", -- $045c1
          17858 => x"80", -- $045c2
          17859 => x"80", -- $045c3
          17860 => x"80", -- $045c4
          17861 => x"7f", -- $045c5
          17862 => x"7f", -- $045c6
          17863 => x"7f", -- $045c7
          17864 => x"7e", -- $045c8
          17865 => x"7e", -- $045c9
          17866 => x"7e", -- $045ca
          17867 => x"7e", -- $045cb
          17868 => x"7e", -- $045cc
          17869 => x"7e", -- $045cd
          17870 => x"7e", -- $045ce
          17871 => x"7e", -- $045cf
          17872 => x"7d", -- $045d0
          17873 => x"7d", -- $045d1
          17874 => x"7d", -- $045d2
          17875 => x"7e", -- $045d3
          17876 => x"7e", -- $045d4
          17877 => x"7f", -- $045d5
          17878 => x"7f", -- $045d6
          17879 => x"80", -- $045d7
          17880 => x"80", -- $045d8
          17881 => x"80", -- $045d9
          17882 => x"80", -- $045da
          17883 => x"81", -- $045db
          17884 => x"81", -- $045dc
          17885 => x"82", -- $045dd
          17886 => x"82", -- $045de
          17887 => x"82", -- $045df
          17888 => x"83", -- $045e0
          17889 => x"83", -- $045e1
          17890 => x"83", -- $045e2
          17891 => x"83", -- $045e3
          17892 => x"83", -- $045e4
          17893 => x"83", -- $045e5
          17894 => x"84", -- $045e6
          17895 => x"84", -- $045e7
          17896 => x"83", -- $045e8
          17897 => x"83", -- $045e9
          17898 => x"83", -- $045ea
          17899 => x"82", -- $045eb
          17900 => x"82", -- $045ec
          17901 => x"81", -- $045ed
          17902 => x"81", -- $045ee
          17903 => x"80", -- $045ef
          17904 => x"80", -- $045f0
          17905 => x"80", -- $045f1
          17906 => x"7f", -- $045f2
          17907 => x"7f", -- $045f3
          17908 => x"7e", -- $045f4
          17909 => x"7e", -- $045f5
          17910 => x"7e", -- $045f6
          17911 => x"7e", -- $045f7
          17912 => x"7e", -- $045f8
          17913 => x"7e", -- $045f9
          17914 => x"7e", -- $045fa
          17915 => x"7e", -- $045fb
          17916 => x"7e", -- $045fc
          17917 => x"7f", -- $045fd
          17918 => x"7f", -- $045fe
          17919 => x"7f", -- $045ff
          17920 => x"7f", -- $04600
          17921 => x"7f", -- $04601
          17922 => x"7f", -- $04602
          17923 => x"7f", -- $04603
          17924 => x"7f", -- $04604
          17925 => x"7f", -- $04605
          17926 => x"7f", -- $04606
          17927 => x"7f", -- $04607
          17928 => x"7f", -- $04608
          17929 => x"80", -- $04609
          17930 => x"80", -- $0460a
          17931 => x"80", -- $0460b
          17932 => x"80", -- $0460c
          17933 => x"80", -- $0460d
          17934 => x"80", -- $0460e
          17935 => x"80", -- $0460f
          17936 => x"80", -- $04610
          17937 => x"80", -- $04611
          17938 => x"80", -- $04612
          17939 => x"80", -- $04613
          17940 => x"80", -- $04614
          17941 => x"80", -- $04615
          17942 => x"80", -- $04616
          17943 => x"80", -- $04617
          17944 => x"80", -- $04618
          17945 => x"80", -- $04619
          17946 => x"80", -- $0461a
          17947 => x"80", -- $0461b
          17948 => x"80", -- $0461c
          17949 => x"80", -- $0461d
          17950 => x"80", -- $0461e
          17951 => x"80", -- $0461f
          17952 => x"80", -- $04620
          17953 => x"80", -- $04621
          17954 => x"80", -- $04622
          17955 => x"80", -- $04623
          17956 => x"80", -- $04624
          17957 => x"80", -- $04625
          17958 => x"80", -- $04626
          17959 => x"81", -- $04627
          17960 => x"81", -- $04628
          17961 => x"81", -- $04629
          17962 => x"81", -- $0462a
          17963 => x"82", -- $0462b
          17964 => x"82", -- $0462c
          17965 => x"82", -- $0462d
          17966 => x"82", -- $0462e
          17967 => x"82", -- $0462f
          17968 => x"82", -- $04630
          17969 => x"82", -- $04631
          17970 => x"82", -- $04632
          17971 => x"81", -- $04633
          17972 => x"81", -- $04634
          17973 => x"80", -- $04635
          17974 => x"80", -- $04636
          17975 => x"80", -- $04637
          17976 => x"80", -- $04638
          17977 => x"80", -- $04639
          17978 => x"80", -- $0463a
          17979 => x"7f", -- $0463b
          17980 => x"7f", -- $0463c
          17981 => x"7f", -- $0463d
          17982 => x"7f", -- $0463e
          17983 => x"7e", -- $0463f
          17984 => x"7e", -- $04640
          17985 => x"7e", -- $04641
          17986 => x"7e", -- $04642
          17987 => x"7e", -- $04643
          17988 => x"7e", -- $04644
          17989 => x"7f", -- $04645
          17990 => x"7f", -- $04646
          17991 => x"7f", -- $04647
          17992 => x"80", -- $04648
          17993 => x"80", -- $04649
          17994 => x"80", -- $0464a
          17995 => x"80", -- $0464b
          17996 => x"80", -- $0464c
          17997 => x"80", -- $0464d
          17998 => x"80", -- $0464e
          17999 => x"81", -- $0464f
          18000 => x"81", -- $04650
          18001 => x"81", -- $04651
          18002 => x"82", -- $04652
          18003 => x"82", -- $04653
          18004 => x"81", -- $04654
          18005 => x"81", -- $04655
          18006 => x"81", -- $04656
          18007 => x"81", -- $04657
          18008 => x"81", -- $04658
          18009 => x"80", -- $04659
          18010 => x"80", -- $0465a
          18011 => x"80", -- $0465b
          18012 => x"80", -- $0465c
          18013 => x"80", -- $0465d
          18014 => x"80", -- $0465e
          18015 => x"80", -- $0465f
          18016 => x"80", -- $04660
          18017 => x"80", -- $04661
          18018 => x"80", -- $04662
          18019 => x"80", -- $04663
          18020 => x"80", -- $04664
          18021 => x"80", -- $04665
          18022 => x"80", -- $04666
          18023 => x"80", -- $04667
          18024 => x"7f", -- $04668
          18025 => x"7f", -- $04669
          18026 => x"7f", -- $0466a
          18027 => x"7f", -- $0466b
          18028 => x"7f", -- $0466c
          18029 => x"7f", -- $0466d
          18030 => x"7f", -- $0466e
          18031 => x"7f", -- $0466f
          18032 => x"7f", -- $04670
          18033 => x"7f", -- $04671
          18034 => x"7f", -- $04672
          18035 => x"7f", -- $04673
          18036 => x"7f", -- $04674
          18037 => x"7f", -- $04675
          18038 => x"7f", -- $04676
          18039 => x"80", -- $04677
          18040 => x"80", -- $04678
          18041 => x"80", -- $04679
          18042 => x"80", -- $0467a
          18043 => x"80", -- $0467b
          18044 => x"80", -- $0467c
          18045 => x"80", -- $0467d
          18046 => x"80", -- $0467e
          18047 => x"80", -- $0467f
          18048 => x"80", -- $04680
          18049 => x"80", -- $04681
          18050 => x"80", -- $04682
          18051 => x"80", -- $04683
          18052 => x"80", -- $04684
          18053 => x"80", -- $04685
          18054 => x"80", -- $04686
          18055 => x"80", -- $04687
          18056 => x"80", -- $04688
          18057 => x"7f", -- $04689
          18058 => x"7f", -- $0468a
          18059 => x"7e", -- $0468b
          18060 => x"7e", -- $0468c
          18061 => x"7e", -- $0468d
          18062 => x"7e", -- $0468e
          18063 => x"7e", -- $0468f
          18064 => x"7e", -- $04690
          18065 => x"7f", -- $04691
          18066 => x"7f", -- $04692
          18067 => x"7f", -- $04693
          18068 => x"80", -- $04694
          18069 => x"80", -- $04695
          18070 => x"80", -- $04696
          18071 => x"80", -- $04697
          18072 => x"80", -- $04698
          18073 => x"80", -- $04699
          18074 => x"80", -- $0469a
          18075 => x"80", -- $0469b
          18076 => x"80", -- $0469c
          18077 => x"80", -- $0469d
          18078 => x"80", -- $0469e
          18079 => x"80", -- $0469f
          18080 => x"81", -- $046a0
          18081 => x"81", -- $046a1
          18082 => x"81", -- $046a2
          18083 => x"81", -- $046a3
          18084 => x"81", -- $046a4
          18085 => x"81", -- $046a5
          18086 => x"81", -- $046a6
          18087 => x"81", -- $046a7
          18088 => x"81", -- $046a8
          18089 => x"80", -- $046a9
          18090 => x"80", -- $046aa
          18091 => x"80", -- $046ab
          18092 => x"80", -- $046ac
          18093 => x"80", -- $046ad
          18094 => x"80", -- $046ae
          18095 => x"80", -- $046af
          18096 => x"80", -- $046b0
          18097 => x"7f", -- $046b1
          18098 => x"7f", -- $046b2
          18099 => x"7f", -- $046b3
          18100 => x"7f", -- $046b4
          18101 => x"7f", -- $046b5
          18102 => x"7f", -- $046b6
          18103 => x"7f", -- $046b7
          18104 => x"7f", -- $046b8
          18105 => x"7f", -- $046b9
          18106 => x"7f", -- $046ba
          18107 => x"7f", -- $046bb
          18108 => x"7f", -- $046bc
          18109 => x"7f", -- $046bd
          18110 => x"7f", -- $046be
          18111 => x"7f", -- $046bf
          18112 => x"7f", -- $046c0
          18113 => x"7f", -- $046c1
          18114 => x"7f", -- $046c2
          18115 => x"80", -- $046c3
          18116 => x"80", -- $046c4
          18117 => x"80", -- $046c5
          18118 => x"80", -- $046c6
          18119 => x"80", -- $046c7
          18120 => x"80", -- $046c8
          18121 => x"80", -- $046c9
          18122 => x"80", -- $046ca
          18123 => x"81", -- $046cb
          18124 => x"81", -- $046cc
          18125 => x"81", -- $046cd
          18126 => x"81", -- $046ce
          18127 => x"80", -- $046cf
          18128 => x"80", -- $046d0
          18129 => x"80", -- $046d1
          18130 => x"80", -- $046d2
          18131 => x"80", -- $046d3
          18132 => x"80", -- $046d4
          18133 => x"80", -- $046d5
          18134 => x"80", -- $046d6
          18135 => x"80", -- $046d7
          18136 => x"80", -- $046d8
          18137 => x"80", -- $046d9
          18138 => x"80", -- $046da
          18139 => x"80", -- $046db
          18140 => x"80", -- $046dc
          18141 => x"80", -- $046dd
          18142 => x"80", -- $046de
          18143 => x"80", -- $046df
          18144 => x"80", -- $046e0
          18145 => x"80", -- $046e1
          18146 => x"80", -- $046e2
          18147 => x"80", -- $046e3
          18148 => x"80", -- $046e4
          18149 => x"80", -- $046e5
          18150 => x"80", -- $046e6
          18151 => x"80", -- $046e7
          18152 => x"80", -- $046e8
          18153 => x"80", -- $046e9
          18154 => x"80", -- $046ea
          18155 => x"80", -- $046eb
          18156 => x"80", -- $046ec
          18157 => x"80", -- $046ed
          18158 => x"80", -- $046ee
          18159 => x"80", -- $046ef
          18160 => x"80", -- $046f0
          18161 => x"80", -- $046f1
          18162 => x"80", -- $046f2
          18163 => x"80", -- $046f3
          18164 => x"80", -- $046f4
          18165 => x"80", -- $046f5
          18166 => x"80", -- $046f6
          18167 => x"80", -- $046f7
          18168 => x"80", -- $046f8
          18169 => x"80", -- $046f9
          18170 => x"80", -- $046fa
          18171 => x"80", -- $046fb
          18172 => x"80", -- $046fc
          18173 => x"80", -- $046fd
          18174 => x"80", -- $046fe
          18175 => x"80", -- $046ff
          18176 => x"80", -- $04700
          18177 => x"80", -- $04701
          18178 => x"80", -- $04702
          18179 => x"80", -- $04703
          18180 => x"80", -- $04704
          18181 => x"7f", -- $04705
          18182 => x"80", -- $04706
          18183 => x"80", -- $04707
          18184 => x"80", -- $04708
          18185 => x"80", -- $04709
          18186 => x"80", -- $0470a
          18187 => x"80", -- $0470b
          18188 => x"80", -- $0470c
          18189 => x"80", -- $0470d
          18190 => x"80", -- $0470e
          18191 => x"80", -- $0470f
          18192 => x"80", -- $04710
          18193 => x"80", -- $04711
          18194 => x"80", -- $04712
          18195 => x"80", -- $04713
          18196 => x"81", -- $04714
          18197 => x"81", -- $04715
          18198 => x"81", -- $04716
          18199 => x"81", -- $04717
          18200 => x"81", -- $04718
          18201 => x"81", -- $04719
          18202 => x"81", -- $0471a
          18203 => x"81", -- $0471b
          18204 => x"81", -- $0471c
          18205 => x"81", -- $0471d
          18206 => x"81", -- $0471e
          18207 => x"81", -- $0471f
          18208 => x"81", -- $04720
          18209 => x"80", -- $04721
          18210 => x"80", -- $04722
          18211 => x"80", -- $04723
          18212 => x"80", -- $04724
          18213 => x"80", -- $04725
          18214 => x"80", -- $04726
          18215 => x"80", -- $04727
          18216 => x"80", -- $04728
          18217 => x"80", -- $04729
          18218 => x"80", -- $0472a
          18219 => x"7f", -- $0472b
          18220 => x"7f", -- $0472c
          18221 => x"7e", -- $0472d
          18222 => x"7c", -- $0472e
          18223 => x"7f", -- $0472f
          18224 => x"80", -- $04730
          18225 => x"80", -- $04731
          18226 => x"7f", -- $04732
          18227 => x"7e", -- $04733
          18228 => x"7f", -- $04734
          18229 => x"7f", -- $04735
          18230 => x"7f", -- $04736
          18231 => x"7f", -- $04737
          18232 => x"80", -- $04738
          18233 => x"7f", -- $04739
          18234 => x"7f", -- $0473a
          18235 => x"80", -- $0473b
          18236 => x"80", -- $0473c
          18237 => x"7f", -- $0473d
          18238 => x"7e", -- $0473e
          18239 => x"7e", -- $0473f
          18240 => x"80", -- $04740
          18241 => x"81", -- $04741
          18242 => x"81", -- $04742
          18243 => x"80", -- $04743
          18244 => x"7f", -- $04744
          18245 => x"7f", -- $04745
          18246 => x"80", -- $04746
          18247 => x"80", -- $04747
          18248 => x"80", -- $04748
          18249 => x"7f", -- $04749
          18250 => x"7f", -- $0474a
          18251 => x"7f", -- $0474b
          18252 => x"7f", -- $0474c
          18253 => x"7f", -- $0474d
          18254 => x"7f", -- $0474e
          18255 => x"80", -- $0474f
          18256 => x"80", -- $04750
          18257 => x"80", -- $04751
          18258 => x"80", -- $04752
          18259 => x"7f", -- $04753
          18260 => x"80", -- $04754
          18261 => x"80", -- $04755
          18262 => x"80", -- $04756
          18263 => x"80", -- $04757
          18264 => x"80", -- $04758
          18265 => x"80", -- $04759
          18266 => x"80", -- $0475a
          18267 => x"7f", -- $0475b
          18268 => x"7f", -- $0475c
          18269 => x"7f", -- $0475d
          18270 => x"80", -- $0475e
          18271 => x"80", -- $0475f
          18272 => x"80", -- $04760
          18273 => x"80", -- $04761
          18274 => x"80", -- $04762
          18275 => x"80", -- $04763
          18276 => x"80", -- $04764
          18277 => x"80", -- $04765
          18278 => x"80", -- $04766
          18279 => x"80", -- $04767
          18280 => x"80", -- $04768
          18281 => x"80", -- $04769
          18282 => x"80", -- $0476a
          18283 => x"80", -- $0476b
          18284 => x"80", -- $0476c
          18285 => x"80", -- $0476d
          18286 => x"80", -- $0476e
          18287 => x"80", -- $0476f
          18288 => x"80", -- $04770
          18289 => x"80", -- $04771
          18290 => x"80", -- $04772
          18291 => x"7f", -- $04773
          18292 => x"7f", -- $04774
          18293 => x"7f", -- $04775
          18294 => x"7f", -- $04776
          18295 => x"7f", -- $04777
          18296 => x"7f", -- $04778
          18297 => x"7f", -- $04779
          18298 => x"7f", -- $0477a
          18299 => x"7f", -- $0477b
          18300 => x"7f", -- $0477c
          18301 => x"7f", -- $0477d
          18302 => x"7f", -- $0477e
          18303 => x"7f", -- $0477f
          18304 => x"80", -- $04780
          18305 => x"80", -- $04781
          18306 => x"80", -- $04782
          18307 => x"80", -- $04783
          18308 => x"80", -- $04784
          18309 => x"80", -- $04785
          18310 => x"80", -- $04786
          18311 => x"80", -- $04787
          18312 => x"80", -- $04788
          18313 => x"80", -- $04789
          18314 => x"80", -- $0478a
          18315 => x"80", -- $0478b
          18316 => x"80", -- $0478c
          18317 => x"80", -- $0478d
          18318 => x"80", -- $0478e
          18319 => x"80", -- $0478f
          18320 => x"80", -- $04790
          18321 => x"80", -- $04791
          18322 => x"80", -- $04792
          18323 => x"80", -- $04793
          18324 => x"80", -- $04794
          18325 => x"80", -- $04795
          18326 => x"80", -- $04796
          18327 => x"80", -- $04797
          18328 => x"80", -- $04798
          18329 => x"80", -- $04799
          18330 => x"80", -- $0479a
          18331 => x"80", -- $0479b
          18332 => x"80", -- $0479c
          18333 => x"80", -- $0479d
          18334 => x"80", -- $0479e
          18335 => x"80", -- $0479f
          18336 => x"80", -- $047a0
          18337 => x"80", -- $047a1
          18338 => x"80", -- $047a2
          18339 => x"80", -- $047a3
          18340 => x"80", -- $047a4
          18341 => x"80", -- $047a5
          18342 => x"80", -- $047a6
          18343 => x"80", -- $047a7
          18344 => x"80", -- $047a8
          18345 => x"80", -- $047a9
          18346 => x"80", -- $047aa
          18347 => x"80", -- $047ab
          18348 => x"80", -- $047ac
          18349 => x"80", -- $047ad
          18350 => x"80", -- $047ae
          18351 => x"80", -- $047af
          18352 => x"80", -- $047b0
          18353 => x"80", -- $047b1
          18354 => x"80", -- $047b2
          18355 => x"80", -- $047b3
          18356 => x"80", -- $047b4
          18357 => x"80", -- $047b5
          18358 => x"80", -- $047b6
          18359 => x"80", -- $047b7
          18360 => x"80", -- $047b8
          18361 => x"80", -- $047b9
          18362 => x"80", -- $047ba
          18363 => x"80", -- $047bb
          18364 => x"80", -- $047bc
          18365 => x"80", -- $047bd
          18366 => x"80", -- $047be
          18367 => x"80", -- $047bf
          18368 => x"80", -- $047c0
          18369 => x"80", -- $047c1
          18370 => x"80", -- $047c2
          18371 => x"80", -- $047c3
          18372 => x"80", -- $047c4
          18373 => x"80", -- $047c5
          18374 => x"80", -- $047c6
          18375 => x"80", -- $047c7
          18376 => x"80", -- $047c8
          18377 => x"80", -- $047c9
          18378 => x"80", -- $047ca
          18379 => x"80", -- $047cb
          18380 => x"80", -- $047cc
          18381 => x"80", -- $047cd
          18382 => x"80", -- $047ce
          18383 => x"80", -- $047cf
          18384 => x"80", -- $047d0
          18385 => x"81", -- $047d1
          18386 => x"80", -- $047d2
          18387 => x"80", -- $047d3
          18388 => x"81", -- $047d4
          18389 => x"80", -- $047d5
          18390 => x"80", -- $047d6
          18391 => x"80", -- $047d7
          18392 => x"80", -- $047d8
          18393 => x"80", -- $047d9
          18394 => x"81", -- $047da
          18395 => x"81", -- $047db
          18396 => x"81", -- $047dc
          18397 => x"81", -- $047dd
          18398 => x"80", -- $047de
          18399 => x"80", -- $047df
          18400 => x"81", -- $047e0
          18401 => x"81", -- $047e1
          18402 => x"81", -- $047e2
          18403 => x"81", -- $047e3
          18404 => x"81", -- $047e4
          18405 => x"80", -- $047e5
          18406 => x"80", -- $047e6
          18407 => x"80", -- $047e7
          18408 => x"80", -- $047e8
          18409 => x"80", -- $047e9
          18410 => x"80", -- $047ea
          18411 => x"80", -- $047eb
          18412 => x"80", -- $047ec
          18413 => x"80", -- $047ed
          18414 => x"80", -- $047ee
          18415 => x"80", -- $047ef
          18416 => x"80", -- $047f0
          18417 => x"80", -- $047f1
          18418 => x"80", -- $047f2
          18419 => x"80", -- $047f3
          18420 => x"80", -- $047f4
          18421 => x"80", -- $047f5
          18422 => x"80", -- $047f6
          18423 => x"80", -- $047f7
          18424 => x"80", -- $047f8
          18425 => x"7f", -- $047f9
          18426 => x"80", -- $047fa
          18427 => x"80", -- $047fb
          18428 => x"80", -- $047fc
          18429 => x"80", -- $047fd
          18430 => x"80", -- $047fe
          18431 => x"80", -- $047ff
          18432 => x"80", -- $04800
          18433 => x"80", -- $04801
          18434 => x"80", -- $04802
          18435 => x"80", -- $04803
          18436 => x"81", -- $04804
          18437 => x"81", -- $04805
          18438 => x"81", -- $04806
          18439 => x"80", -- $04807
          18440 => x"80", -- $04808
          18441 => x"80", -- $04809
          18442 => x"80", -- $0480a
          18443 => x"80", -- $0480b
          18444 => x"80", -- $0480c
          18445 => x"80", -- $0480d
          18446 => x"80", -- $0480e
          18447 => x"80", -- $0480f
          18448 => x"80", -- $04810
          18449 => x"80", -- $04811
          18450 => x"80", -- $04812
          18451 => x"80", -- $04813
          18452 => x"80", -- $04814
          18453 => x"80", -- $04815
          18454 => x"80", -- $04816
          18455 => x"80", -- $04817
          18456 => x"80", -- $04818
          18457 => x"80", -- $04819
          18458 => x"80", -- $0481a
          18459 => x"80", -- $0481b
          18460 => x"80", -- $0481c
          18461 => x"80", -- $0481d
          18462 => x"80", -- $0481e
          18463 => x"80", -- $0481f
          18464 => x"80", -- $04820
          18465 => x"80", -- $04821
          18466 => x"81", -- $04822
          18467 => x"81", -- $04823
          18468 => x"80", -- $04824
          18469 => x"80", -- $04825
          18470 => x"80", -- $04826
          18471 => x"80", -- $04827
          18472 => x"80", -- $04828
          18473 => x"80", -- $04829
          18474 => x"80", -- $0482a
          18475 => x"80", -- $0482b
          18476 => x"80", -- $0482c
          18477 => x"80", -- $0482d
          18478 => x"7f", -- $0482e
          18479 => x"7f", -- $0482f
          18480 => x"7f", -- $04830
          18481 => x"7f", -- $04831
          18482 => x"80", -- $04832
          18483 => x"80", -- $04833
          18484 => x"80", -- $04834
          18485 => x"80", -- $04835
          18486 => x"80", -- $04836
          18487 => x"80", -- $04837
          18488 => x"80", -- $04838
          18489 => x"80", -- $04839
          18490 => x"80", -- $0483a
          18491 => x"80", -- $0483b
          18492 => x"80", -- $0483c
          18493 => x"80", -- $0483d
          18494 => x"80", -- $0483e
          18495 => x"80", -- $0483f
          18496 => x"80", -- $04840
          18497 => x"80", -- $04841
          18498 => x"80", -- $04842
          18499 => x"80", -- $04843
          18500 => x"80", -- $04844
          18501 => x"80", -- $04845
          18502 => x"80", -- $04846
          18503 => x"80", -- $04847
          18504 => x"80", -- $04848
          18505 => x"80", -- $04849
          18506 => x"80", -- $0484a
          18507 => x"80", -- $0484b
          18508 => x"80", -- $0484c
          18509 => x"80", -- $0484d
          18510 => x"80", -- $0484e
          18511 => x"80", -- $0484f
          18512 => x"80", -- $04850
          18513 => x"80", -- $04851
          18514 => x"80", -- $04852
          18515 => x"80", -- $04853
          18516 => x"80", -- $04854
          18517 => x"80", -- $04855
          18518 => x"80", -- $04856
          18519 => x"80", -- $04857
          18520 => x"80", -- $04858
          18521 => x"80", -- $04859
          18522 => x"80", -- $0485a
          18523 => x"80", -- $0485b
          18524 => x"80", -- $0485c
          18525 => x"80", -- $0485d
          18526 => x"80", -- $0485e
          18527 => x"80", -- $0485f
          18528 => x"80", -- $04860
          18529 => x"80", -- $04861
          18530 => x"80", -- $04862
          18531 => x"80", -- $04863
          18532 => x"80", -- $04864
          18533 => x"80", -- $04865
          18534 => x"80", -- $04866
          18535 => x"80", -- $04867
          18536 => x"80", -- $04868
          18537 => x"80", -- $04869
          18538 => x"80", -- $0486a
          18539 => x"80", -- $0486b
          18540 => x"80", -- $0486c
          18541 => x"80", -- $0486d
          18542 => x"80", -- $0486e
          18543 => x"80", -- $0486f
          18544 => x"80", -- $04870
          18545 => x"80", -- $04871
          18546 => x"80", -- $04872
          18547 => x"80", -- $04873
          18548 => x"81", -- $04874
          18549 => x"81", -- $04875
          18550 => x"81", -- $04876
          18551 => x"81", -- $04877
          18552 => x"80", -- $04878
          18553 => x"80", -- $04879
          18554 => x"80", -- $0487a
          18555 => x"80", -- $0487b
          18556 => x"80", -- $0487c
          18557 => x"80", -- $0487d
          18558 => x"80", -- $0487e
          18559 => x"80", -- $0487f
          18560 => x"81", -- $04880
          18561 => x"81", -- $04881
          18562 => x"80", -- $04882
          18563 => x"80", -- $04883
          18564 => x"80", -- $04884
          18565 => x"80", -- $04885
          18566 => x"81", -- $04886
          18567 => x"81", -- $04887
          18568 => x"81", -- $04888
          18569 => x"81", -- $04889
          18570 => x"80", -- $0488a
          18571 => x"80", -- $0488b
          18572 => x"80", -- $0488c
          18573 => x"80", -- $0488d
          18574 => x"80", -- $0488e
          18575 => x"80", -- $0488f
          18576 => x"80", -- $04890
          18577 => x"80", -- $04891
          18578 => x"81", -- $04892
          18579 => x"81", -- $04893
          18580 => x"81", -- $04894
          18581 => x"80", -- $04895
          18582 => x"80", -- $04896
          18583 => x"80", -- $04897
          18584 => x"80", -- $04898
          18585 => x"80", -- $04899
          18586 => x"80", -- $0489a
          18587 => x"80", -- $0489b
          18588 => x"80", -- $0489c
          18589 => x"80", -- $0489d
          18590 => x"80", -- $0489e
          18591 => x"80", -- $0489f
          18592 => x"80", -- $048a0
          18593 => x"80", -- $048a1
          18594 => x"7f", -- $048a2
          18595 => x"7f", -- $048a3
          18596 => x"7f", -- $048a4
          18597 => x"7f", -- $048a5
          18598 => x"7f", -- $048a6
          18599 => x"7f", -- $048a7
          18600 => x"7f", -- $048a8
          18601 => x"7f", -- $048a9
          18602 => x"7f", -- $048aa
          18603 => x"7f", -- $048ab
          18604 => x"7f", -- $048ac
          18605 => x"7f", -- $048ad
          18606 => x"7f", -- $048ae
          18607 => x"7f", -- $048af
          18608 => x"7f", -- $048b0
          18609 => x"7f", -- $048b1
          18610 => x"80", -- $048b2
          18611 => x"80", -- $048b3
          18612 => x"80", -- $048b4
          18613 => x"80", -- $048b5
          18614 => x"81", -- $048b6
          18615 => x"81", -- $048b7
          18616 => x"82", -- $048b8
          18617 => x"83", -- $048b9
          18618 => x"84", -- $048ba
          18619 => x"85", -- $048bb
          18620 => x"84", -- $048bc
          18621 => x"84", -- $048bd
          18622 => x"83", -- $048be
          18623 => x"83", -- $048bf
          18624 => x"83", -- $048c0
          18625 => x"84", -- $048c1
          18626 => x"84", -- $048c2
          18627 => x"85", -- $048c3
          18628 => x"85", -- $048c4
          18629 => x"84", -- $048c5
          18630 => x"83", -- $048c6
          18631 => x"82", -- $048c7
          18632 => x"81", -- $048c8
          18633 => x"81", -- $048c9
          18634 => x"81", -- $048ca
          18635 => x"81", -- $048cb
          18636 => x"80", -- $048cc
          18637 => x"80", -- $048cd
          18638 => x"7e", -- $048ce
          18639 => x"7e", -- $048cf
          18640 => x"7e", -- $048d0
          18641 => x"7f", -- $048d1
          18642 => x"7f", -- $048d2
          18643 => x"7f", -- $048d3
          18644 => x"7e", -- $048d4
          18645 => x"7c", -- $048d5
          18646 => x"7a", -- $048d6
          18647 => x"7a", -- $048d7
          18648 => x"7a", -- $048d8
          18649 => x"7c", -- $048d9
          18650 => x"7d", -- $048da
          18651 => x"7e", -- $048db
          18652 => x"7e", -- $048dc
          18653 => x"7e", -- $048dd
          18654 => x"7c", -- $048de
          18655 => x"7c", -- $048df
          18656 => x"7c", -- $048e0
          18657 => x"7c", -- $048e1
          18658 => x"7c", -- $048e2
          18659 => x"7d", -- $048e3
          18660 => x"7c", -- $048e4
          18661 => x"7c", -- $048e5
          18662 => x"7d", -- $048e6
          18663 => x"7d", -- $048e7
          18664 => x"7f", -- $048e8
          18665 => x"80", -- $048e9
          18666 => x"81", -- $048ea
          18667 => x"81", -- $048eb
          18668 => x"81", -- $048ec
          18669 => x"81", -- $048ed
          18670 => x"81", -- $048ee
          18671 => x"83", -- $048ef
          18672 => x"85", -- $048f0
          18673 => x"85", -- $048f1
          18674 => x"87", -- $048f2
          18675 => x"86", -- $048f3
          18676 => x"86", -- $048f4
          18677 => x"86", -- $048f5
          18678 => x"86", -- $048f6
          18679 => x"88", -- $048f7
          18680 => x"89", -- $048f8
          18681 => x"88", -- $048f9
          18682 => x"86", -- $048fa
          18683 => x"82", -- $048fb
          18684 => x"80", -- $048fc
          18685 => x"7e", -- $048fd
          18686 => x"80", -- $048fe
          18687 => x"80", -- $048ff
          18688 => x"84", -- $04900
          18689 => x"85", -- $04901
          18690 => x"84", -- $04902
          18691 => x"81", -- $04903
          18692 => x"7e", -- $04904
          18693 => x"7b", -- $04905
          18694 => x"79", -- $04906
          18695 => x"79", -- $04907
          18696 => x"7a", -- $04908
          18697 => x"7a", -- $04909
          18698 => x"7b", -- $0490a
          18699 => x"7a", -- $0490b
          18700 => x"7b", -- $0490c
          18701 => x"7c", -- $0490d
          18702 => x"7e", -- $0490e
          18703 => x"81", -- $0490f
          18704 => x"84", -- $04910
          18705 => x"86", -- $04911
          18706 => x"86", -- $04912
          18707 => x"85", -- $04913
          18708 => x"81", -- $04914
          18709 => x"80", -- $04915
          18710 => x"7f", -- $04916
          18711 => x"7e", -- $04917
          18712 => x"7e", -- $04918
          18713 => x"7c", -- $04919
          18714 => x"7a", -- $0491a
          18715 => x"76", -- $0491b
          18716 => x"75", -- $0491c
          18717 => x"74", -- $0491d
          18718 => x"75", -- $0491e
          18719 => x"77", -- $0491f
          18720 => x"7a", -- $04920
          18721 => x"7d", -- $04921
          18722 => x"7e", -- $04922
          18723 => x"7f", -- $04923
          18724 => x"80", -- $04924
          18725 => x"80", -- $04925
          18726 => x"81", -- $04926
          18727 => x"82", -- $04927
          18728 => x"82", -- $04928
          18729 => x"81", -- $04929
          18730 => x"80", -- $0492a
          18731 => x"7e", -- $0492b
          18732 => x"7c", -- $0492c
          18733 => x"7c", -- $0492d
          18734 => x"7d", -- $0492e
          18735 => x"7f", -- $0492f
          18736 => x"81", -- $04930
          18737 => x"82", -- $04931
          18738 => x"84", -- $04932
          18739 => x"85", -- $04933
          18740 => x"85", -- $04934
          18741 => x"87", -- $04935
          18742 => x"87", -- $04936
          18743 => x"88", -- $04937
          18744 => x"88", -- $04938
          18745 => x"87", -- $04939
          18746 => x"86", -- $0493a
          18747 => x"84", -- $0493b
          18748 => x"83", -- $0493c
          18749 => x"83", -- $0493d
          18750 => x"84", -- $0493e
          18751 => x"86", -- $0493f
          18752 => x"84", -- $04940
          18753 => x"82", -- $04941
          18754 => x"81", -- $04942
          18755 => x"80", -- $04943
          18756 => x"80", -- $04944
          18757 => x"81", -- $04945
          18758 => x"83", -- $04946
          18759 => x"85", -- $04947
          18760 => x"84", -- $04948
          18761 => x"83", -- $04949
          18762 => x"80", -- $0494a
          18763 => x"7d", -- $0494b
          18764 => x"7a", -- $0494c
          18765 => x"79", -- $0494d
          18766 => x"7a", -- $0494e
          18767 => x"7a", -- $0494f
          18768 => x"7c", -- $04950
          18769 => x"7b", -- $04951
          18770 => x"7b", -- $04952
          18771 => x"7b", -- $04953
          18772 => x"7a", -- $04954
          18773 => x"7c", -- $04955
          18774 => x"7f", -- $04956
          18775 => x"80", -- $04957
          18776 => x"81", -- $04958
          18777 => x"81", -- $04959
          18778 => x"80", -- $0495a
          18779 => x"7f", -- $0495b
          18780 => x"7c", -- $0495c
          18781 => x"7a", -- $0495d
          18782 => x"78", -- $0495e
          18783 => x"77", -- $0495f
          18784 => x"77", -- $04960
          18785 => x"77", -- $04961
          18786 => x"78", -- $04962
          18787 => x"78", -- $04963
          18788 => x"7a", -- $04964
          18789 => x"7d", -- $04965
          18790 => x"7f", -- $04966
          18791 => x"81", -- $04967
          18792 => x"83", -- $04968
          18793 => x"84", -- $04969
          18794 => x"85", -- $0496a
          18795 => x"85", -- $0496b
          18796 => x"84", -- $0496c
          18797 => x"84", -- $0496d
          18798 => x"83", -- $0496e
          18799 => x"82", -- $0496f
          18800 => x"82", -- $04970
          18801 => x"81", -- $04971
          18802 => x"80", -- $04972
          18803 => x"80", -- $04973
          18804 => x"80", -- $04974
          18805 => x"81", -- $04975
          18806 => x"83", -- $04976
          18807 => x"86", -- $04977
          18808 => x"8a", -- $04978
          18809 => x"8c", -- $04979
          18810 => x"8c", -- $0497a
          18811 => x"8c", -- $0497b
          18812 => x"8b", -- $0497c
          18813 => x"88", -- $0497d
          18814 => x"87", -- $0497e
          18815 => x"86", -- $0497f
          18816 => x"85", -- $04980
          18817 => x"85", -- $04981
          18818 => x"83", -- $04982
          18819 => x"82", -- $04983
          18820 => x"80", -- $04984
          18821 => x"7e", -- $04985
          18822 => x"7c", -- $04986
          18823 => x"7b", -- $04987
          18824 => x"7a", -- $04988
          18825 => x"7c", -- $04989
          18826 => x"7d", -- $0498a
          18827 => x"7e", -- $0498b
          18828 => x"7f", -- $0498c
          18829 => x"80", -- $0498d
          18830 => x"80", -- $0498e
          18831 => x"80", -- $0498f
          18832 => x"80", -- $04990
          18833 => x"80", -- $04991
          18834 => x"80", -- $04992
          18835 => x"81", -- $04993
          18836 => x"81", -- $04994
          18837 => x"81", -- $04995
          18838 => x"80", -- $04996
          18839 => x"80", -- $04997
          18840 => x"7f", -- $04998
          18841 => x"7e", -- $04999
          18842 => x"7c", -- $0499a
          18843 => x"7b", -- $0499b
          18844 => x"79", -- $0499c
          18845 => x"78", -- $0499d
          18846 => x"76", -- $0499e
          18847 => x"75", -- $0499f
          18848 => x"74", -- $049a0
          18849 => x"73", -- $049a1
          18850 => x"74", -- $049a2
          18851 => x"74", -- $049a3
          18852 => x"76", -- $049a4
          18853 => x"79", -- $049a5
          18854 => x"7b", -- $049a6
          18855 => x"7e", -- $049a7
          18856 => x"80", -- $049a8
          18857 => x"82", -- $049a9
          18858 => x"84", -- $049aa
          18859 => x"86", -- $049ab
          18860 => x"87", -- $049ac
          18861 => x"88", -- $049ad
          18862 => x"88", -- $049ae
          18863 => x"87", -- $049af
          18864 => x"86", -- $049b0
          18865 => x"85", -- $049b1
          18866 => x"84", -- $049b2
          18867 => x"83", -- $049b3
          18868 => x"82", -- $049b4
          18869 => x"81", -- $049b5
          18870 => x"81", -- $049b6
          18871 => x"81", -- $049b7
          18872 => x"82", -- $049b8
          18873 => x"83", -- $049b9
          18874 => x"84", -- $049ba
          18875 => x"86", -- $049bb
          18876 => x"87", -- $049bc
          18877 => x"88", -- $049bd
          18878 => x"89", -- $049be
          18879 => x"89", -- $049bf
          18880 => x"89", -- $049c0
          18881 => x"88", -- $049c1
          18882 => x"87", -- $049c2
          18883 => x"86", -- $049c3
          18884 => x"85", -- $049c4
          18885 => x"84", -- $049c5
          18886 => x"82", -- $049c6
          18887 => x"80", -- $049c7
          18888 => x"7f", -- $049c8
          18889 => x"7d", -- $049c9
          18890 => x"7e", -- $049ca
          18891 => x"7d", -- $049cb
          18892 => x"7f", -- $049cc
          18893 => x"7f", -- $049cd
          18894 => x"80", -- $049ce
          18895 => x"80", -- $049cf
          18896 => x"80", -- $049d0
          18897 => x"7e", -- $049d1
          18898 => x"7c", -- $049d2
          18899 => x"7c", -- $049d3
          18900 => x"7a", -- $049d4
          18901 => x"7b", -- $049d5
          18902 => x"79", -- $049d6
          18903 => x"79", -- $049d7
          18904 => x"77", -- $049d8
          18905 => x"76", -- $049d9
          18906 => x"76", -- $049da
          18907 => x"75", -- $049db
          18908 => x"77", -- $049dc
          18909 => x"78", -- $049dd
          18910 => x"7a", -- $049de
          18911 => x"7b", -- $049df
          18912 => x"7c", -- $049e0
          18913 => x"7d", -- $049e1
          18914 => x"7e", -- $049e2
          18915 => x"7f", -- $049e3
          18916 => x"7f", -- $049e4
          18917 => x"80", -- $049e5
          18918 => x"80", -- $049e6
          18919 => x"80", -- $049e7
          18920 => x"7f", -- $049e8
          18921 => x"7f", -- $049e9
          18922 => x"7e", -- $049ea
          18923 => x"7e", -- $049eb
          18924 => x"7f", -- $049ec
          18925 => x"7f", -- $049ed
          18926 => x"80", -- $049ee
          18927 => x"80", -- $049ef
          18928 => x"80", -- $049f0
          18929 => x"81", -- $049f1
          18930 => x"82", -- $049f2
          18931 => x"83", -- $049f3
          18932 => x"85", -- $049f4
          18933 => x"86", -- $049f5
          18934 => x"86", -- $049f6
          18935 => x"87", -- $049f7
          18936 => x"87", -- $049f8
          18937 => x"87", -- $049f9
          18938 => x"87", -- $049fa
          18939 => x"88", -- $049fb
          18940 => x"88", -- $049fc
          18941 => x"89", -- $049fd
          18942 => x"8a", -- $049fe
          18943 => x"8a", -- $049ff
          18944 => x"89", -- $04a00
          18945 => x"88", -- $04a01
          18946 => x"87", -- $04a02
          18947 => x"87", -- $04a03
          18948 => x"85", -- $04a04
          18949 => x"86", -- $04a05
          18950 => x"85", -- $04a06
          18951 => x"84", -- $04a07
          18952 => x"83", -- $04a08
          18953 => x"80", -- $04a09
          18954 => x"7f", -- $04a0a
          18955 => x"7c", -- $04a0b
          18956 => x"7b", -- $04a0c
          18957 => x"79", -- $04a0d
          18958 => x"79", -- $04a0e
          18959 => x"78", -- $04a0f
          18960 => x"78", -- $04a10
          18961 => x"78", -- $04a11
          18962 => x"77", -- $04a12
          18963 => x"77", -- $04a13
          18964 => x"78", -- $04a14
          18965 => x"79", -- $04a15
          18966 => x"7a", -- $04a16
          18967 => x"7c", -- $04a17
          18968 => x"7e", -- $04a18
          18969 => x"7f", -- $04a19
          18970 => x"80", -- $04a1a
          18971 => x"80", -- $04a1b
          18972 => x"80", -- $04a1c
          18973 => x"80", -- $04a1d
          18974 => x"80", -- $04a1e
          18975 => x"80", -- $04a1f
          18976 => x"80", -- $04a20
          18977 => x"7f", -- $04a21
          18978 => x"7d", -- $04a22
          18979 => x"7c", -- $04a23
          18980 => x"7a", -- $04a24
          18981 => x"79", -- $04a25
          18982 => x"79", -- $04a26
          18983 => x"78", -- $04a27
          18984 => x"79", -- $04a28
          18985 => x"78", -- $04a29
          18986 => x"79", -- $04a2a
          18987 => x"7a", -- $04a2b
          18988 => x"7c", -- $04a2c
          18989 => x"7e", -- $04a2d
          18990 => x"80", -- $04a2e
          18991 => x"82", -- $04a2f
          18992 => x"84", -- $04a30
          18993 => x"86", -- $04a31
          18994 => x"87", -- $04a32
          18995 => x"88", -- $04a33
          18996 => x"88", -- $04a34
          18997 => x"89", -- $04a35
          18998 => x"88", -- $04a36
          18999 => x"89", -- $04a37
          19000 => x"88", -- $04a38
          19001 => x"87", -- $04a39
          19002 => x"86", -- $04a3a
          19003 => x"84", -- $04a3b
          19004 => x"83", -- $04a3c
          19005 => x"82", -- $04a3d
          19006 => x"81", -- $04a3e
          19007 => x"80", -- $04a3f
          19008 => x"81", -- $04a40
          19009 => x"81", -- $04a41
          19010 => x"81", -- $04a42
          19011 => x"82", -- $04a43
          19012 => x"82", -- $04a44
          19013 => x"83", -- $04a45
          19014 => x"84", -- $04a46
          19015 => x"85", -- $04a47
          19016 => x"85", -- $04a48
          19017 => x"86", -- $04a49
          19018 => x"85", -- $04a4a
          19019 => x"86", -- $04a4b
          19020 => x"85", -- $04a4c
          19021 => x"83", -- $04a4d
          19022 => x"82", -- $04a4e
          19023 => x"80", -- $04a4f
          19024 => x"80", -- $04a50
          19025 => x"7e", -- $04a51
          19026 => x"7c", -- $04a52
          19027 => x"7d", -- $04a53
          19028 => x"7a", -- $04a54
          19029 => x"7a", -- $04a55
          19030 => x"79", -- $04a56
          19031 => x"78", -- $04a57
          19032 => x"78", -- $04a58
          19033 => x"78", -- $04a59
          19034 => x"78", -- $04a5a
          19035 => x"79", -- $04a5b
          19036 => x"79", -- $04a5c
          19037 => x"79", -- $04a5d
          19038 => x"7a", -- $04a5e
          19039 => x"79", -- $04a5f
          19040 => x"7b", -- $04a60
          19041 => x"7b", -- $04a61
          19042 => x"7c", -- $04a62
          19043 => x"7c", -- $04a63
          19044 => x"7c", -- $04a64
          19045 => x"7e", -- $04a65
          19046 => x"7d", -- $04a66
          19047 => x"7e", -- $04a67
          19048 => x"7e", -- $04a68
          19049 => x"7f", -- $04a69
          19050 => x"7f", -- $04a6a
          19051 => x"7f", -- $04a6b
          19052 => x"7f", -- $04a6c
          19053 => x"7f", -- $04a6d
          19054 => x"80", -- $04a6e
          19055 => x"7f", -- $04a6f
          19056 => x"80", -- $04a70
          19057 => x"80", -- $04a71
          19058 => x"80", -- $04a72
          19059 => x"81", -- $04a73
          19060 => x"81", -- $04a74
          19061 => x"81", -- $04a75
          19062 => x"82", -- $04a76
          19063 => x"82", -- $04a77
          19064 => x"83", -- $04a78
          19065 => x"84", -- $04a79
          19066 => x"85", -- $04a7a
          19067 => x"85", -- $04a7b
          19068 => x"86", -- $04a7c
          19069 => x"85", -- $04a7d
          19070 => x"86", -- $04a7e
          19071 => x"85", -- $04a7f
          19072 => x"85", -- $04a80
          19073 => x"85", -- $04a81
          19074 => x"85", -- $04a82
          19075 => x"85", -- $04a83
          19076 => x"85", -- $04a84
          19077 => x"85", -- $04a85
          19078 => x"85", -- $04a86
          19079 => x"84", -- $04a87
          19080 => x"84", -- $04a88
          19081 => x"83", -- $04a89
          19082 => x"82", -- $04a8a
          19083 => x"82", -- $04a8b
          19084 => x"81", -- $04a8c
          19085 => x"81", -- $04a8d
          19086 => x"80", -- $04a8e
          19087 => x"80", -- $04a8f
          19088 => x"7f", -- $04a90
          19089 => x"7d", -- $04a91
          19090 => x"7c", -- $04a92
          19091 => x"7b", -- $04a93
          19092 => x"7a", -- $04a94
          19093 => x"79", -- $04a95
          19094 => x"79", -- $04a96
          19095 => x"78", -- $04a97
          19096 => x"78", -- $04a98
          19097 => x"77", -- $04a99
          19098 => x"78", -- $04a9a
          19099 => x"78", -- $04a9b
          19100 => x"79", -- $04a9c
          19101 => x"7a", -- $04a9d
          19102 => x"7c", -- $04a9e
          19103 => x"7e", -- $04a9f
          19104 => x"7f", -- $04aa0
          19105 => x"80", -- $04aa1
          19106 => x"80", -- $04aa2
          19107 => x"80", -- $04aa3
          19108 => x"81", -- $04aa4
          19109 => x"81", -- $04aa5
          19110 => x"81", -- $04aa6
          19111 => x"80", -- $04aa7
          19112 => x"80", -- $04aa8
          19113 => x"7f", -- $04aa9
          19114 => x"7d", -- $04aaa
          19115 => x"7c", -- $04aab
          19116 => x"7b", -- $04aac
          19117 => x"7a", -- $04aad
          19118 => x"7a", -- $04aae
          19119 => x"7a", -- $04aaf
          19120 => x"7a", -- $04ab0
          19121 => x"7a", -- $04ab1
          19122 => x"7b", -- $04ab2
          19123 => x"7c", -- $04ab3
          19124 => x"7e", -- $04ab4
          19125 => x"7f", -- $04ab5
          19126 => x"80", -- $04ab6
          19127 => x"82", -- $04ab7
          19128 => x"83", -- $04ab8
          19129 => x"84", -- $04ab9
          19130 => x"85", -- $04aba
          19131 => x"85", -- $04abb
          19132 => x"86", -- $04abc
          19133 => x"86", -- $04abd
          19134 => x"86", -- $04abe
          19135 => x"86", -- $04abf
          19136 => x"85", -- $04ac0
          19137 => x"83", -- $04ac1
          19138 => x"83", -- $04ac2
          19139 => x"82", -- $04ac3
          19140 => x"81", -- $04ac4
          19141 => x"81", -- $04ac5
          19142 => x"80", -- $04ac6
          19143 => x"80", -- $04ac7
          19144 => x"80", -- $04ac8
          19145 => x"80", -- $04ac9
          19146 => x"7f", -- $04aca
          19147 => x"80", -- $04acb
          19148 => x"80", -- $04acc
          19149 => x"81", -- $04acd
          19150 => x"82", -- $04ace
          19151 => x"82", -- $04acf
          19152 => x"82", -- $04ad0
          19153 => x"82", -- $04ad1
          19154 => x"82", -- $04ad2
          19155 => x"82", -- $04ad3
          19156 => x"82", -- $04ad4
          19157 => x"81", -- $04ad5
          19158 => x"81", -- $04ad6
          19159 => x"80", -- $04ad7
          19160 => x"7f", -- $04ad8
          19161 => x"7f", -- $04ad9
          19162 => x"7c", -- $04ada
          19163 => x"7d", -- $04adb
          19164 => x"7d", -- $04adc
          19165 => x"7c", -- $04add
          19166 => x"7e", -- $04ade
          19167 => x"7c", -- $04adf
          19168 => x"7d", -- $04ae0
          19169 => x"7d", -- $04ae1
          19170 => x"7d", -- $04ae2
          19171 => x"7d", -- $04ae3
          19172 => x"7f", -- $04ae4
          19173 => x"7f", -- $04ae5
          19174 => x"7f", -- $04ae6
          19175 => x"80", -- $04ae7
          19176 => x"7e", -- $04ae8
          19177 => x"7f", -- $04ae9
          19178 => x"7e", -- $04aea
          19179 => x"7f", -- $04aeb
          19180 => x"7f", -- $04aec
          19181 => x"80", -- $04aed
          19182 => x"7f", -- $04aee
          19183 => x"7e", -- $04aef
          19184 => x"7e", -- $04af0
          19185 => x"7e", -- $04af1
          19186 => x"7f", -- $04af2
          19187 => x"80", -- $04af3
          19188 => x"80", -- $04af4
          19189 => x"80", -- $04af5
          19190 => x"81", -- $04af6
          19191 => x"80", -- $04af7
          19192 => x"80", -- $04af8
          19193 => x"80", -- $04af9
          19194 => x"80", -- $04afa
          19195 => x"81", -- $04afb
          19196 => x"81", -- $04afc
          19197 => x"81", -- $04afd
          19198 => x"80", -- $04afe
          19199 => x"80", -- $04aff
          19200 => x"80", -- $04b00
          19201 => x"80", -- $04b01
          19202 => x"81", -- $04b02
          19203 => x"82", -- $04b03
          19204 => x"82", -- $04b04
          19205 => x"83", -- $04b05
          19206 => x"83", -- $04b06
          19207 => x"82", -- $04b07
          19208 => x"83", -- $04b08
          19209 => x"83", -- $04b09
          19210 => x"84", -- $04b0a
          19211 => x"84", -- $04b0b
          19212 => x"85", -- $04b0c
          19213 => x"85", -- $04b0d
          19214 => x"84", -- $04b0e
          19215 => x"84", -- $04b0f
          19216 => x"85", -- $04b10
          19217 => x"84", -- $04b11
          19218 => x"84", -- $04b12
          19219 => x"84", -- $04b13
          19220 => x"82", -- $04b14
          19221 => x"83", -- $04b15
          19222 => x"81", -- $04b16
          19223 => x"81", -- $04b17
          19224 => x"81", -- $04b18
          19225 => x"80", -- $04b19
          19226 => x"80", -- $04b1a
          19227 => x"80", -- $04b1b
          19228 => x"7f", -- $04b1c
          19229 => x"7d", -- $04b1d
          19230 => x"7d", -- $04b1e
          19231 => x"7c", -- $04b1f
          19232 => x"7c", -- $04b20
          19233 => x"7b", -- $04b21
          19234 => x"7b", -- $04b22
          19235 => x"7a", -- $04b23
          19236 => x"7a", -- $04b24
          19237 => x"7b", -- $04b25
          19238 => x"7b", -- $04b26
          19239 => x"7c", -- $04b27
          19240 => x"7d", -- $04b28
          19241 => x"7e", -- $04b29
          19242 => x"7f", -- $04b2a
          19243 => x"80", -- $04b2b
          19244 => x"80", -- $04b2c
          19245 => x"82", -- $04b2d
          19246 => x"82", -- $04b2e
          19247 => x"83", -- $04b2f
          19248 => x"83", -- $04b30
          19249 => x"82", -- $04b31
          19250 => x"82", -- $04b32
          19251 => x"82", -- $04b33
          19252 => x"82", -- $04b34
          19253 => x"81", -- $04b35
          19254 => x"80", -- $04b36
          19255 => x"80", -- $04b37
          19256 => x"7f", -- $04b38
          19257 => x"7f", -- $04b39
          19258 => x"7e", -- $04b3a
          19259 => x"7e", -- $04b3b
          19260 => x"7e", -- $04b3c
          19261 => x"7e", -- $04b3d
          19262 => x"7e", -- $04b3e
          19263 => x"7e", -- $04b3f
          19264 => x"7f", -- $04b40
          19265 => x"7f", -- $04b41
          19266 => x"80", -- $04b42
          19267 => x"80", -- $04b43
          19268 => x"80", -- $04b44
          19269 => x"80", -- $04b45
          19270 => x"81", -- $04b46
          19271 => x"81", -- $04b47
          19272 => x"81", -- $04b48
          19273 => x"82", -- $04b49
          19274 => x"82", -- $04b4a
          19275 => x"83", -- $04b4b
          19276 => x"83", -- $04b4c
          19277 => x"82", -- $04b4d
          19278 => x"82", -- $04b4e
          19279 => x"82", -- $04b4f
          19280 => x"82", -- $04b50
          19281 => x"82", -- $04b51
          19282 => x"81", -- $04b52
          19283 => x"81", -- $04b53
          19284 => x"81", -- $04b54
          19285 => x"81", -- $04b55
          19286 => x"81", -- $04b56
          19287 => x"81", -- $04b57
          19288 => x"81", -- $04b58
          19289 => x"81", -- $04b59
          19290 => x"81", -- $04b5a
          19291 => x"81", -- $04b5b
          19292 => x"80", -- $04b5c
          19293 => x"81", -- $04b5d
          19294 => x"81", -- $04b5e
          19295 => x"81", -- $04b5f
          19296 => x"81", -- $04b60
          19297 => x"80", -- $04b61
          19298 => x"80", -- $04b62
          19299 => x"80", -- $04b63
          19300 => x"80", -- $04b64
          19301 => x"80", -- $04b65
          19302 => x"80", -- $04b66
          19303 => x"7f", -- $04b67
          19304 => x"7e", -- $04b68
          19305 => x"80", -- $04b69
          19306 => x"7f", -- $04b6a
          19307 => x"80", -- $04b6b
          19308 => x"80", -- $04b6c
          19309 => x"81", -- $04b6d
          19310 => x"81", -- $04b6e
          19311 => x"80", -- $04b6f
          19312 => x"80", -- $04b70
          19313 => x"80", -- $04b71
          19314 => x"81", -- $04b72
          19315 => x"81", -- $04b73
          19316 => x"80", -- $04b74
          19317 => x"80", -- $04b75
          19318 => x"7f", -- $04b76
          19319 => x"7e", -- $04b77
          19320 => x"7e", -- $04b78
          19321 => x"7d", -- $04b79
          19322 => x"7d", -- $04b7a
          19323 => x"7b", -- $04b7b
          19324 => x"7b", -- $04b7c
          19325 => x"7b", -- $04b7d
          19326 => x"7c", -- $04b7e
          19327 => x"7d", -- $04b7f
          19328 => x"7d", -- $04b80
          19329 => x"7e", -- $04b81
          19330 => x"7e", -- $04b82
          19331 => x"7f", -- $04b83
          19332 => x"80", -- $04b84
          19333 => x"80", -- $04b85
          19334 => x"81", -- $04b86
          19335 => x"80", -- $04b87
          19336 => x"80", -- $04b88
          19337 => x"80", -- $04b89
          19338 => x"80", -- $04b8a
          19339 => x"80", -- $04b8b
          19340 => x"80", -- $04b8c
          19341 => x"7f", -- $04b8d
          19342 => x"7f", -- $04b8e
          19343 => x"80", -- $04b8f
          19344 => x"80", -- $04b90
          19345 => x"81", -- $04b91
          19346 => x"80", -- $04b92
          19347 => x"80", -- $04b93
          19348 => x"82", -- $04b94
          19349 => x"84", -- $04b95
          19350 => x"85", -- $04b96
          19351 => x"85", -- $04b97
          19352 => x"85", -- $04b98
          19353 => x"86", -- $04b99
          19354 => x"88", -- $04b9a
          19355 => x"88", -- $04b9b
          19356 => x"87", -- $04b9c
          19357 => x"82", -- $04b9d
          19358 => x"82", -- $04b9e
          19359 => x"81", -- $04b9f
          19360 => x"82", -- $04ba0
          19361 => x"84", -- $04ba1
          19362 => x"81", -- $04ba2
          19363 => x"81", -- $04ba3
          19364 => x"80", -- $04ba4
          19365 => x"82", -- $04ba5
          19366 => x"82", -- $04ba6
          19367 => x"81", -- $04ba7
          19368 => x"80", -- $04ba8
          19369 => x"7d", -- $04ba9
          19370 => x"7e", -- $04baa
          19371 => x"7d", -- $04bab
          19372 => x"7c", -- $04bac
          19373 => x"7b", -- $04bad
          19374 => x"79", -- $04bae
          19375 => x"7a", -- $04baf
          19376 => x"7c", -- $04bb0
          19377 => x"7e", -- $04bb1
          19378 => x"7f", -- $04bb2
          19379 => x"7f", -- $04bb3
          19380 => x"80", -- $04bb4
          19381 => x"83", -- $04bb5
          19382 => x"85", -- $04bb6
          19383 => x"85", -- $04bb7
          19384 => x"84", -- $04bb8
          19385 => x"84", -- $04bb9
          19386 => x"83", -- $04bba
          19387 => x"82", -- $04bbb
          19388 => x"80", -- $04bbc
          19389 => x"7d", -- $04bbd
          19390 => x"7a", -- $04bbe
          19391 => x"79", -- $04bbf
          19392 => x"78", -- $04bc0
          19393 => x"78", -- $04bc1
          19394 => x"79", -- $04bc2
          19395 => x"79", -- $04bc3
          19396 => x"7b", -- $04bc4
          19397 => x"7d", -- $04bc5
          19398 => x"80", -- $04bc6
          19399 => x"81", -- $04bc7
          19400 => x"83", -- $04bc8
          19401 => x"84", -- $04bc9
          19402 => x"84", -- $04bca
          19403 => x"85", -- $04bcb
          19404 => x"83", -- $04bcc
          19405 => x"82", -- $04bcd
          19406 => x"81", -- $04bce
          19407 => x"7f", -- $04bcf
          19408 => x"7d", -- $04bd0
          19409 => x"7c", -- $04bd1
          19410 => x"7b", -- $04bd2
          19411 => x"7b", -- $04bd3
          19412 => x"7b", -- $04bd4
          19413 => x"7c", -- $04bd5
          19414 => x"7e", -- $04bd6
          19415 => x"80", -- $04bd7
          19416 => x"82", -- $04bd8
          19417 => x"84", -- $04bd9
          19418 => x"86", -- $04bda
          19419 => x"86", -- $04bdb
          19420 => x"87", -- $04bdc
          19421 => x"87", -- $04bdd
          19422 => x"85", -- $04bde
          19423 => x"84", -- $04bdf
          19424 => x"82", -- $04be0
          19425 => x"82", -- $04be1
          19426 => x"80", -- $04be2
          19427 => x"80", -- $04be3
          19428 => x"7f", -- $04be4
          19429 => x"7e", -- $04be5
          19430 => x"7f", -- $04be6
          19431 => x"80", -- $04be7
          19432 => x"80", -- $04be8
          19433 => x"80", -- $04be9
          19434 => x"82", -- $04bea
          19435 => x"82", -- $04beb
          19436 => x"82", -- $04bec
          19437 => x"83", -- $04bed
          19438 => x"84", -- $04bee
          19439 => x"83", -- $04bef
          19440 => x"83", -- $04bf0
          19441 => x"82", -- $04bf1
          19442 => x"83", -- $04bf2
          19443 => x"82", -- $04bf3
          19444 => x"80", -- $04bf4
          19445 => x"7e", -- $04bf5
          19446 => x"80", -- $04bf6
          19447 => x"80", -- $04bf7
          19448 => x"80", -- $04bf8
          19449 => x"80", -- $04bf9
          19450 => x"80", -- $04bfa
          19451 => x"81", -- $04bfb
          19452 => x"81", -- $04bfc
          19453 => x"80", -- $04bfd
          19454 => x"80", -- $04bfe
          19455 => x"80", -- $04bff
          19456 => x"7f", -- $04c00
          19457 => x"7e", -- $04c01
          19458 => x"7c", -- $04c02
          19459 => x"7a", -- $04c03
          19460 => x"7b", -- $04c04
          19461 => x"7b", -- $04c05
          19462 => x"7b", -- $04c06
          19463 => x"7b", -- $04c07
          19464 => x"7d", -- $04c08
          19465 => x"80", -- $04c09
          19466 => x"80", -- $04c0a
          19467 => x"81", -- $04c0b
          19468 => x"82", -- $04c0c
          19469 => x"83", -- $04c0d
          19470 => x"85", -- $04c0e
          19471 => x"83", -- $04c0f
          19472 => x"82", -- $04c10
          19473 => x"7f", -- $04c11
          19474 => x"7e", -- $04c12
          19475 => x"7f", -- $04c13
          19476 => x"7b", -- $04c14
          19477 => x"7a", -- $04c15
          19478 => x"78", -- $04c16
          19479 => x"7b", -- $04c17
          19480 => x"7b", -- $04c18
          19481 => x"7b", -- $04c19
          19482 => x"7c", -- $04c1a
          19483 => x"7f", -- $04c1b
          19484 => x"82", -- $04c1c
          19485 => x"83", -- $04c1d
          19486 => x"85", -- $04c1e
          19487 => x"86", -- $04c1f
          19488 => x"89", -- $04c20
          19489 => x"8a", -- $04c21
          19490 => x"88", -- $04c22
          19491 => x"88", -- $04c23
          19492 => x"89", -- $04c24
          19493 => x"87", -- $04c25
          19494 => x"85", -- $04c26
          19495 => x"84", -- $04c27
          19496 => x"84", -- $04c28
          19497 => x"84", -- $04c29
          19498 => x"85", -- $04c2a
          19499 => x"84", -- $04c2b
          19500 => x"80", -- $04c2c
          19501 => x"84", -- $04c2d
          19502 => x"86", -- $04c2e
          19503 => x"85", -- $04c2f
          19504 => x"85", -- $04c30
          19505 => x"84", -- $04c31
          19506 => x"87", -- $04c32
          19507 => x"86", -- $04c33
          19508 => x"83", -- $04c34
          19509 => x"82", -- $04c35
          19510 => x"80", -- $04c36
          19511 => x"7f", -- $04c37
          19512 => x"7c", -- $04c38
          19513 => x"79", -- $04c39
          19514 => x"78", -- $04c3a
          19515 => x"78", -- $04c3b
          19516 => x"77", -- $04c3c
          19517 => x"76", -- $04c3d
          19518 => x"78", -- $04c3e
          19519 => x"7a", -- $04c3f
          19520 => x"7c", -- $04c40
          19521 => x"7e", -- $04c41
          19522 => x"7f", -- $04c42
          19523 => x"81", -- $04c43
          19524 => x"83", -- $04c44
          19525 => x"84", -- $04c45
          19526 => x"84", -- $04c46
          19527 => x"84", -- $04c47
          19528 => x"84", -- $04c48
          19529 => x"82", -- $04c49
          19530 => x"80", -- $04c4a
          19531 => x"7f", -- $04c4b
          19532 => x"7d", -- $04c4c
          19533 => x"7b", -- $04c4d
          19534 => x"7a", -- $04c4e
          19535 => x"79", -- $04c4f
          19536 => x"78", -- $04c50
          19537 => x"79", -- $04c51
          19538 => x"7a", -- $04c52
          19539 => x"7a", -- $04c53
          19540 => x"7c", -- $04c54
          19541 => x"7d", -- $04c55
          19542 => x"7f", -- $04c56
          19543 => x"80", -- $04c57
          19544 => x"80", -- $04c58
          19545 => x"80", -- $04c59
          19546 => x"81", -- $04c5a
          19547 => x"82", -- $04c5b
          19548 => x"80", -- $04c5c
          19549 => x"80", -- $04c5d
          19550 => x"80", -- $04c5e
          19551 => x"80", -- $04c5f
          19552 => x"7f", -- $04c60
          19553 => x"7e", -- $04c61
          19554 => x"7e", -- $04c62
          19555 => x"7f", -- $04c63
          19556 => x"80", -- $04c64
          19557 => x"7f", -- $04c65
          19558 => x"80", -- $04c66
          19559 => x"80", -- $04c67
          19560 => x"81", -- $04c68
          19561 => x"81", -- $04c69
          19562 => x"81", -- $04c6a
          19563 => x"83", -- $04c6b
          19564 => x"83", -- $04c6c
          19565 => x"82", -- $04c6d
          19566 => x"82", -- $04c6e
          19567 => x"83", -- $04c6f
          19568 => x"83", -- $04c70
          19569 => x"82", -- $04c71
          19570 => x"82", -- $04c72
          19571 => x"82", -- $04c73
          19572 => x"83", -- $04c74
          19573 => x"82", -- $04c75
          19574 => x"82", -- $04c76
          19575 => x"82", -- $04c77
          19576 => x"80", -- $04c78
          19577 => x"81", -- $04c79
          19578 => x"80", -- $04c7a
          19579 => x"80", -- $04c7b
          19580 => x"80", -- $04c7c
          19581 => x"7f", -- $04c7d
          19582 => x"7f", -- $04c7e
          19583 => x"80", -- $04c7f
          19584 => x"80", -- $04c80
          19585 => x"81", -- $04c81
          19586 => x"81", -- $04c82
          19587 => x"80", -- $04c83
          19588 => x"81", -- $04c84
          19589 => x"83", -- $04c85
          19590 => x"83", -- $04c86
          19591 => x"82", -- $04c87
          19592 => x"82", -- $04c88
          19593 => x"83", -- $04c89
          19594 => x"82", -- $04c8a
          19595 => x"80", -- $04c8b
          19596 => x"80", -- $04c8c
          19597 => x"80", -- $04c8d
          19598 => x"7e", -- $04c8e
          19599 => x"7c", -- $04c8f
          19600 => x"7b", -- $04c90
          19601 => x"7b", -- $04c91
          19602 => x"7b", -- $04c92
          19603 => x"7a", -- $04c93
          19604 => x"7a", -- $04c94
          19605 => x"7d", -- $04c95
          19606 => x"7e", -- $04c96
          19607 => x"80", -- $04c97
          19608 => x"80", -- $04c98
          19609 => x"81", -- $04c99
          19610 => x"83", -- $04c9a
          19611 => x"83", -- $04c9b
          19612 => x"82", -- $04c9c
          19613 => x"83", -- $04c9d
          19614 => x"82", -- $04c9e
          19615 => x"80", -- $04c9f
          19616 => x"80", -- $04ca0
          19617 => x"7e", -- $04ca1
          19618 => x"7e", -- $04ca2
          19619 => x"7c", -- $04ca3
          19620 => x"7b", -- $04ca4
          19621 => x"7b", -- $04ca5
          19622 => x"7b", -- $04ca6
          19623 => x"7c", -- $04ca7
          19624 => x"7d", -- $04ca8
          19625 => x"7f", -- $04ca9
          19626 => x"80", -- $04caa
          19627 => x"81", -- $04cab
          19628 => x"83", -- $04cac
          19629 => x"84", -- $04cad
          19630 => x"86", -- $04cae
          19631 => x"87", -- $04caf
          19632 => x"88", -- $04cb0
          19633 => x"88", -- $04cb1
          19634 => x"88", -- $04cb2
          19635 => x"87", -- $04cb3
          19636 => x"85", -- $04cb4
          19637 => x"87", -- $04cb5
          19638 => x"86", -- $04cb6
          19639 => x"85", -- $04cb7
          19640 => x"84", -- $04cb8
          19641 => x"82", -- $04cb9
          19642 => x"81", -- $04cba
          19643 => x"83", -- $04cbb
          19644 => x"81", -- $04cbc
          19645 => x"81", -- $04cbd
          19646 => x"82", -- $04cbe
          19647 => x"83", -- $04cbf
          19648 => x"83", -- $04cc0
          19649 => x"81", -- $04cc1
          19650 => x"82", -- $04cc2
          19651 => x"83", -- $04cc3
          19652 => x"81", -- $04cc4
          19653 => x"80", -- $04cc5
          19654 => x"7f", -- $04cc6
          19655 => x"7e", -- $04cc7
          19656 => x"7d", -- $04cc8
          19657 => x"7b", -- $04cc9
          19658 => x"7a", -- $04cca
          19659 => x"7a", -- $04ccb
          19660 => x"7b", -- $04ccc
          19661 => x"7a", -- $04ccd
          19662 => x"7b", -- $04cce
          19663 => x"7d", -- $04ccf
          19664 => x"7e", -- $04cd0
          19665 => x"7f", -- $04cd1
          19666 => x"80", -- $04cd2
          19667 => x"81", -- $04cd3
          19668 => x"82", -- $04cd4
          19669 => x"83", -- $04cd5
          19670 => x"83", -- $04cd6
          19671 => x"83", -- $04cd7
          19672 => x"83", -- $04cd8
          19673 => x"81", -- $04cd9
          19674 => x"80", -- $04cda
          19675 => x"80", -- $04cdb
          19676 => x"7f", -- $04cdc
          19677 => x"7d", -- $04cdd
          19678 => x"7c", -- $04cde
          19679 => x"7b", -- $04cdf
          19680 => x"7b", -- $04ce0
          19681 => x"7a", -- $04ce1
          19682 => x"7b", -- $04ce2
          19683 => x"7b", -- $04ce3
          19684 => x"7c", -- $04ce4
          19685 => x"7e", -- $04ce5
          19686 => x"7f", -- $04ce6
          19687 => x"80", -- $04ce7
          19688 => x"80", -- $04ce8
          19689 => x"81", -- $04ce9
          19690 => x"81", -- $04cea
          19691 => x"81", -- $04ceb
          19692 => x"82", -- $04cec
          19693 => x"82", -- $04ced
          19694 => x"82", -- $04cee
          19695 => x"82", -- $04cef
          19696 => x"81", -- $04cf0
          19697 => x"80", -- $04cf1
          19698 => x"80", -- $04cf2
          19699 => x"80", -- $04cf3
          19700 => x"80", -- $04cf4
          19701 => x"80", -- $04cf5
          19702 => x"7f", -- $04cf6
          19703 => x"80", -- $04cf7
          19704 => x"7f", -- $04cf8
          19705 => x"7f", -- $04cf9
          19706 => x"80", -- $04cfa
          19707 => x"7f", -- $04cfb
          19708 => x"80", -- $04cfc
          19709 => x"80", -- $04cfd
          19710 => x"81", -- $04cfe
          19711 => x"80", -- $04cff
          19712 => x"82", -- $04d00
          19713 => x"82", -- $04d01
          19714 => x"82", -- $04d02
          19715 => x"82", -- $04d03
          19716 => x"82", -- $04d04
          19717 => x"83", -- $04d05
          19718 => x"81", -- $04d06
          19719 => x"80", -- $04d07
          19720 => x"80", -- $04d08
          19721 => x"80", -- $04d09
          19722 => x"7e", -- $04d0a
          19723 => x"7d", -- $04d0b
          19724 => x"7d", -- $04d0c
          19725 => x"7d", -- $04d0d
          19726 => x"7c", -- $04d0e
          19727 => x"7d", -- $04d0f
          19728 => x"7e", -- $04d10
          19729 => x"7e", -- $04d11
          19730 => x"7f", -- $04d12
          19731 => x"80", -- $04d13
          19732 => x"80", -- $04d14
          19733 => x"82", -- $04d15
          19734 => x"82", -- $04d16
          19735 => x"82", -- $04d17
          19736 => x"82", -- $04d18
          19737 => x"82", -- $04d19
          19738 => x"81", -- $04d1a
          19739 => x"80", -- $04d1b
          19740 => x"80", -- $04d1c
          19741 => x"7f", -- $04d1d
          19742 => x"7d", -- $04d1e
          19743 => x"7c", -- $04d1f
          19744 => x"7c", -- $04d20
          19745 => x"7b", -- $04d21
          19746 => x"7b", -- $04d22
          19747 => x"7b", -- $04d23
          19748 => x"7c", -- $04d24
          19749 => x"7c", -- $04d25
          19750 => x"7e", -- $04d26
          19751 => x"7f", -- $04d27
          19752 => x"80", -- $04d28
          19753 => x"80", -- $04d29
          19754 => x"81", -- $04d2a
          19755 => x"81", -- $04d2b
          19756 => x"81", -- $04d2c
          19757 => x"81", -- $04d2d
          19758 => x"80", -- $04d2e
          19759 => x"80", -- $04d2f
          19760 => x"7f", -- $04d30
          19761 => x"7f", -- $04d31
          19762 => x"7e", -- $04d32
          19763 => x"7e", -- $04d33
          19764 => x"7d", -- $04d34
          19765 => x"7e", -- $04d35
          19766 => x"7e", -- $04d36
          19767 => x"7f", -- $04d37
          19768 => x"80", -- $04d38
          19769 => x"80", -- $04d39
          19770 => x"81", -- $04d3a
          19771 => x"82", -- $04d3b
          19772 => x"83", -- $04d3c
          19773 => x"84", -- $04d3d
          19774 => x"86", -- $04d3e
          19775 => x"86", -- $04d3f
          19776 => x"87", -- $04d40
          19777 => x"88", -- $04d41
          19778 => x"86", -- $04d42
          19779 => x"85", -- $04d43
          19780 => x"86", -- $04d44
          19781 => x"83", -- $04d45
          19782 => x"82", -- $04d46
          19783 => x"82", -- $04d47
          19784 => x"81", -- $04d48
          19785 => x"80", -- $04d49
          19786 => x"7f", -- $04d4a
          19787 => x"7f", -- $04d4b
          19788 => x"7f", -- $04d4c
          19789 => x"7d", -- $04d4d
          19790 => x"7d", -- $04d4e
          19791 => x"7d", -- $04d4f
          19792 => x"7c", -- $04d50
          19793 => x"7b", -- $04d51
          19794 => x"7b", -- $04d52
          19795 => x"7c", -- $04d53
          19796 => x"7b", -- $04d54
          19797 => x"7b", -- $04d55
          19798 => x"7c", -- $04d56
          19799 => x"7d", -- $04d57
          19800 => x"7e", -- $04d58
          19801 => x"7f", -- $04d59
          19802 => x"80", -- $04d5a
          19803 => x"80", -- $04d5b
          19804 => x"81", -- $04d5c
          19805 => x"81", -- $04d5d
          19806 => x"82", -- $04d5e
          19807 => x"82", -- $04d5f
          19808 => x"82", -- $04d60
          19809 => x"81", -- $04d61
          19810 => x"80", -- $04d62
          19811 => x"80", -- $04d63
          19812 => x"7e", -- $04d64
          19813 => x"7d", -- $04d65
          19814 => x"7c", -- $04d66
          19815 => x"7a", -- $04d67
          19816 => x"7a", -- $04d68
          19817 => x"7a", -- $04d69
          19818 => x"79", -- $04d6a
          19819 => x"7a", -- $04d6b
          19820 => x"7a", -- $04d6c
          19821 => x"7c", -- $04d6d
          19822 => x"7d", -- $04d6e
          19823 => x"7d", -- $04d6f
          19824 => x"7f", -- $04d70
          19825 => x"80", -- $04d71
          19826 => x"80", -- $04d72
          19827 => x"80", -- $04d73
          19828 => x"80", -- $04d74
          19829 => x"82", -- $04d75
          19830 => x"80", -- $04d76
          19831 => x"80", -- $04d77
          19832 => x"80", -- $04d78
          19833 => x"80", -- $04d79
          19834 => x"7e", -- $04d7a
          19835 => x"7e", -- $04d7b
          19836 => x"7f", -- $04d7c
          19837 => x"7e", -- $04d7d
          19838 => x"7e", -- $04d7e
          19839 => x"7e", -- $04d7f
          19840 => x"80", -- $04d80
          19841 => x"80", -- $04d81
          19842 => x"80", -- $04d82
          19843 => x"80", -- $04d83
          19844 => x"81", -- $04d84
          19845 => x"81", -- $04d85
          19846 => x"81", -- $04d86
          19847 => x"82", -- $04d87
          19848 => x"82", -- $04d88
          19849 => x"81", -- $04d89
          19850 => x"81", -- $04d8a
          19851 => x"82", -- $04d8b
          19852 => x"82", -- $04d8c
          19853 => x"81", -- $04d8d
          19854 => x"80", -- $04d8e
          19855 => x"80", -- $04d8f
          19856 => x"80", -- $04d90
          19857 => x"7f", -- $04d91
          19858 => x"7e", -- $04d92
          19859 => x"7f", -- $04d93
          19860 => x"7d", -- $04d94
          19861 => x"7d", -- $04d95
          19862 => x"7d", -- $04d96
          19863 => x"7d", -- $04d97
          19864 => x"7d", -- $04d98
          19865 => x"7d", -- $04d99
          19866 => x"7e", -- $04d9a
          19867 => x"7f", -- $04d9b
          19868 => x"7f", -- $04d9c
          19869 => x"80", -- $04d9d
          19870 => x"80", -- $04d9e
          19871 => x"81", -- $04d9f
          19872 => x"81", -- $04da0
          19873 => x"81", -- $04da1
          19874 => x"82", -- $04da2
          19875 => x"81", -- $04da3
          19876 => x"81", -- $04da4
          19877 => x"80", -- $04da5
          19878 => x"80", -- $04da6
          19879 => x"80", -- $04da7
          19880 => x"7f", -- $04da8
          19881 => x"7f", -- $04da9
          19882 => x"7e", -- $04daa
          19883 => x"7e", -- $04dab
          19884 => x"7d", -- $04dac
          19885 => x"7d", -- $04dad
          19886 => x"7d", -- $04dae
          19887 => x"7d", -- $04daf
          19888 => x"7d", -- $04db0
          19889 => x"7e", -- $04db1
          19890 => x"7e", -- $04db2
          19891 => x"7f", -- $04db3
          19892 => x"7f", -- $04db4
          19893 => x"7f", -- $04db5
          19894 => x"80", -- $04db6
          19895 => x"80", -- $04db7
          19896 => x"7f", -- $04db8
          19897 => x"80", -- $04db9
          19898 => x"80", -- $04dba
          19899 => x"80", -- $04dbb
          19900 => x"80", -- $04dbc
          19901 => x"80", -- $04dbd
          19902 => x"80", -- $04dbe
          19903 => x"80", -- $04dbf
          19904 => x"81", -- $04dc0
          19905 => x"83", -- $04dc1
          19906 => x"84", -- $04dc2
          19907 => x"85", -- $04dc3
          19908 => x"86", -- $04dc4
          19909 => x"87", -- $04dc5
          19910 => x"86", -- $04dc6
          19911 => x"88", -- $04dc7
          19912 => x"85", -- $04dc8
          19913 => x"85", -- $04dc9
          19914 => x"87", -- $04dca
          19915 => x"83", -- $04dcb
          19916 => x"83", -- $04dcc
          19917 => x"82", -- $04dcd
          19918 => x"80", -- $04dce
          19919 => x"80", -- $04dcf
          19920 => x"7e", -- $04dd0
          19921 => x"7e", -- $04dd1
          19922 => x"7d", -- $04dd2
          19923 => x"7b", -- $04dd3
          19924 => x"7a", -- $04dd4
          19925 => x"7a", -- $04dd5
          19926 => x"7a", -- $04dd6
          19927 => x"79", -- $04dd7
          19928 => x"7a", -- $04dd8
          19929 => x"7b", -- $04dd9
          19930 => x"7c", -- $04dda
          19931 => x"7c", -- $04ddb
          19932 => x"7e", -- $04ddc
          19933 => x"80", -- $04ddd
          19934 => x"80", -- $04dde
          19935 => x"81", -- $04ddf
          19936 => x"82", -- $04de0
          19937 => x"83", -- $04de1
          19938 => x"83", -- $04de2
          19939 => x"83", -- $04de3
          19940 => x"84", -- $04de4
          19941 => x"83", -- $04de5
          19942 => x"81", -- $04de6
          19943 => x"81", -- $04de7
          19944 => x"80", -- $04de8
          19945 => x"7f", -- $04de9
          19946 => x"7d", -- $04dea
          19947 => x"7c", -- $04deb
          19948 => x"7b", -- $04dec
          19949 => x"79", -- $04ded
          19950 => x"79", -- $04dee
          19951 => x"79", -- $04def
          19952 => x"78", -- $04df0
          19953 => x"79", -- $04df1
          19954 => x"7a", -- $04df2
          19955 => x"7b", -- $04df3
          19956 => x"7c", -- $04df4
          19957 => x"7e", -- $04df5
          19958 => x"7f", -- $04df6
          19959 => x"80", -- $04df7
          19960 => x"80", -- $04df8
          19961 => x"81", -- $04df9
          19962 => x"81", -- $04dfa
          19963 => x"80", -- $04dfb
          19964 => x"82", -- $04dfc
          19965 => x"81", -- $04dfd
          19966 => x"80", -- $04dfe
          19967 => x"80", -- $04dff
          19968 => x"80", -- $04e00
          19969 => x"80", -- $04e01
          19970 => x"7e", -- $04e02
          19971 => x"7e", -- $04e03
          19972 => x"7e", -- $04e04
          19973 => x"7e", -- $04e05
          19974 => x"7d", -- $04e06
          19975 => x"7e", -- $04e07
          19976 => x"7e", -- $04e08
          19977 => x"7e", -- $04e09
          19978 => x"7e", -- $04e0a
          19979 => x"80", -- $04e0b
          19980 => x"80", -- $04e0c
          19981 => x"80", -- $04e0d
          19982 => x"81", -- $04e0e
          19983 => x"81", -- $04e0f
          19984 => x"83", -- $04e10
          19985 => x"82", -- $04e11
          19986 => x"83", -- $04e12
          19987 => x"83", -- $04e13
          19988 => x"83", -- $04e14
          19989 => x"83", -- $04e15
          19990 => x"82", -- $04e16
          19991 => x"81", -- $04e17
          19992 => x"80", -- $04e18
          19993 => x"80", -- $04e19
          19994 => x"7f", -- $04e1a
          19995 => x"7e", -- $04e1b
          19996 => x"7e", -- $04e1c
          19997 => x"7d", -- $04e1d
          19998 => x"7d", -- $04e1e
          19999 => x"7d", -- $04e1f
          20000 => x"7c", -- $04e20
          20001 => x"7d", -- $04e21
          20002 => x"7d", -- $04e22
          20003 => x"7d", -- $04e23
          20004 => x"7e", -- $04e24
          20005 => x"7e", -- $04e25
          20006 => x"7f", -- $04e26
          20007 => x"7f", -- $04e27
          20008 => x"80", -- $04e28
          20009 => x"80", -- $04e29
          20010 => x"80", -- $04e2a
          20011 => x"80", -- $04e2b
          20012 => x"80", -- $04e2c
          20013 => x"80", -- $04e2d
          20014 => x"80", -- $04e2e
          20015 => x"80", -- $04e2f
          20016 => x"80", -- $04e30
          20017 => x"7f", -- $04e31
          20018 => x"7f", -- $04e32
          20019 => x"7f", -- $04e33
          20020 => x"7f", -- $04e34
          20021 => x"80", -- $04e35
          20022 => x"80", -- $04e36
          20023 => x"80", -- $04e37
          20024 => x"80", -- $04e38
          20025 => x"80", -- $04e39
          20026 => x"80", -- $04e3a
          20027 => x"80", -- $04e3b
          20028 => x"80", -- $04e3c
          20029 => x"80", -- $04e3d
          20030 => x"80", -- $04e3e
          20031 => x"80", -- $04e3f
          20032 => x"80", -- $04e40
          20033 => x"80", -- $04e41
          20034 => x"7f", -- $04e42
          20035 => x"80", -- $04e43
          20036 => x"80", -- $04e44
          20037 => x"80", -- $04e45
          20038 => x"80", -- $04e46
          20039 => x"81", -- $04e47
          20040 => x"82", -- $04e48
          20041 => x"82", -- $04e49
          20042 => x"83", -- $04e4a
          20043 => x"85", -- $04e4b
          20044 => x"85", -- $04e4c
          20045 => x"86", -- $04e4d
          20046 => x"86", -- $04e4e
          20047 => x"85", -- $04e4f
          20048 => x"87", -- $04e50
          20049 => x"85", -- $04e51
          20050 => x"85", -- $04e52
          20051 => x"85", -- $04e53
          20052 => x"84", -- $04e54
          20053 => x"83", -- $04e55
          20054 => x"82", -- $04e56
          20055 => x"82", -- $04e57
          20056 => x"80", -- $04e58
          20057 => x"80", -- $04e59
          20058 => x"7f", -- $04e5a
          20059 => x"7f", -- $04e5b
          20060 => x"7d", -- $04e5c
          20061 => x"7d", -- $04e5d
          20062 => x"7d", -- $04e5e
          20063 => x"7d", -- $04e5f
          20064 => x"7c", -- $04e60
          20065 => x"7d", -- $04e61
          20066 => x"7d", -- $04e62
          20067 => x"7e", -- $04e63
          20068 => x"7e", -- $04e64
          20069 => x"7f", -- $04e65
          20070 => x"80", -- $04e66
          20071 => x"80", -- $04e67
          20072 => x"81", -- $04e68
          20073 => x"82", -- $04e69
          20074 => x"83", -- $04e6a
          20075 => x"83", -- $04e6b
          20076 => x"83", -- $04e6c
          20077 => x"83", -- $04e6d
          20078 => x"83", -- $04e6e
          20079 => x"82", -- $04e6f
          20080 => x"82", -- $04e70
          20081 => x"80", -- $04e71
          20082 => x"80", -- $04e72
          20083 => x"7f", -- $04e73
          20084 => x"7e", -- $04e74
          20085 => x"7e", -- $04e75
          20086 => x"7c", -- $04e76
          20087 => x"7d", -- $04e77
          20088 => x"7d", -- $04e78
          20089 => x"7d", -- $04e79
          20090 => x"7e", -- $04e7a
          20091 => x"7e", -- $04e7b
          20092 => x"7f", -- $04e7c
          20093 => x"80", -- $04e7d
          20094 => x"80", -- $04e7e
          20095 => x"80", -- $04e7f
          20096 => x"82", -- $04e80
          20097 => x"82", -- $04e81
          20098 => x"81", -- $04e82
          20099 => x"82", -- $04e83
          20100 => x"83", -- $04e84
          20101 => x"82", -- $04e85
          20102 => x"81", -- $04e86
          20103 => x"82", -- $04e87
          20104 => x"82", -- $04e88
          20105 => x"81", -- $04e89
          20106 => x"80", -- $04e8a
          20107 => x"82", -- $04e8b
          20108 => x"81", -- $04e8c
          20109 => x"80", -- $04e8d
          20110 => x"81", -- $04e8e
          20111 => x"82", -- $04e8f
          20112 => x"82", -- $04e90
          20113 => x"80", -- $04e91
          20114 => x"82", -- $04e92
          20115 => x"83", -- $04e93
          20116 => x"82", -- $04e94
          20117 => x"83", -- $04e95
          20118 => x"84", -- $04e96
          20119 => x"84", -- $04e97
          20120 => x"83", -- $04e98
          20121 => x"84", -- $04e99
          20122 => x"84", -- $04e9a
          20123 => x"83", -- $04e9b
          20124 => x"83", -- $04e9c
          20125 => x"83", -- $04e9d
          20126 => x"82", -- $04e9e
          20127 => x"81", -- $04e9f
          20128 => x"80", -- $04ea0
          20129 => x"80", -- $04ea1
          20130 => x"80", -- $04ea2
          20131 => x"7f", -- $04ea3
          20132 => x"80", -- $04ea4
          20133 => x"7f", -- $04ea5
          20134 => x"7e", -- $04ea6
          20135 => x"7e", -- $04ea7
          20136 => x"80", -- $04ea8
          20137 => x"80", -- $04ea9
          20138 => x"80", -- $04eaa
          20139 => x"80", -- $04eab
          20140 => x"81", -- $04eac
          20141 => x"81", -- $04ead
          20142 => x"81", -- $04eae
          20143 => x"82", -- $04eaf
          20144 => x"82", -- $04eb0
          20145 => x"81", -- $04eb1
          20146 => x"81", -- $04eb2
          20147 => x"81", -- $04eb3
          20148 => x"81", -- $04eb4
          20149 => x"80", -- $04eb5
          20150 => x"80", -- $04eb6
          20151 => x"80", -- $04eb7
          20152 => x"80", -- $04eb8
          20153 => x"7f", -- $04eb9
          20154 => x"7f", -- $04eba
          20155 => x"7f", -- $04ebb
          20156 => x"7f", -- $04ebc
          20157 => x"7f", -- $04ebd
          20158 => x"80", -- $04ebe
          20159 => x"80", -- $04ebf
          20160 => x"80", -- $04ec0
          20161 => x"80", -- $04ec1
          20162 => x"80", -- $04ec2
          20163 => x"80", -- $04ec3
          20164 => x"80", -- $04ec4
          20165 => x"80", -- $04ec5
          20166 => x"80", -- $04ec6
          20167 => x"80", -- $04ec7
          20168 => x"80", -- $04ec8
          20169 => x"80", -- $04ec9
          20170 => x"81", -- $04eca
          20171 => x"81", -- $04ecb
          20172 => x"81", -- $04ecc
          20173 => x"82", -- $04ecd
          20174 => x"83", -- $04ece
          20175 => x"83", -- $04ecf
          20176 => x"84", -- $04ed0
          20177 => x"85", -- $04ed1
          20178 => x"86", -- $04ed2
          20179 => x"86", -- $04ed3
          20180 => x"87", -- $04ed4
          20181 => x"87", -- $04ed5
          20182 => x"87", -- $04ed6
          20183 => x"88", -- $04ed7
          20184 => x"87", -- $04ed8
          20185 => x"86", -- $04ed9
          20186 => x"86", -- $04eda
          20187 => x"85", -- $04edb
          20188 => x"84", -- $04edc
          20189 => x"82", -- $04edd
          20190 => x"82", -- $04ede
          20191 => x"81", -- $04edf
          20192 => x"80", -- $04ee0
          20193 => x"7f", -- $04ee1
          20194 => x"7f", -- $04ee2
          20195 => x"7d", -- $04ee3
          20196 => x"7c", -- $04ee4
          20197 => x"7d", -- $04ee5
          20198 => x"7c", -- $04ee6
          20199 => x"7c", -- $04ee7
          20200 => x"7c", -- $04ee8
          20201 => x"7d", -- $04ee9
          20202 => x"7d", -- $04eea
          20203 => x"7d", -- $04eeb
          20204 => x"7e", -- $04eec
          20205 => x"7f", -- $04eed
          20206 => x"80", -- $04eee
          20207 => x"80", -- $04eef
          20208 => x"81", -- $04ef0
          20209 => x"82", -- $04ef1
          20210 => x"83", -- $04ef2
          20211 => x"83", -- $04ef3
          20212 => x"84", -- $04ef4
          20213 => x"84", -- $04ef5
          20214 => x"84", -- $04ef6
          20215 => x"83", -- $04ef7
          20216 => x"82", -- $04ef8
          20217 => x"81", -- $04ef9
          20218 => x"80", -- $04efa
          20219 => x"80", -- $04efb
          20220 => x"7e", -- $04efc
          20221 => x"7e", -- $04efd
          20222 => x"7e", -- $04efe
          20223 => x"7c", -- $04eff
          20224 => x"7d", -- $04f00
          20225 => x"7d", -- $04f01
          20226 => x"7d", -- $04f02
          20227 => x"7d", -- $04f03
          20228 => x"7e", -- $04f04
          20229 => x"80", -- $04f05
          20230 => x"7e", -- $04f06
          20231 => x"80", -- $04f07
          20232 => x"80", -- $04f08
          20233 => x"81", -- $04f09
          20234 => x"80", -- $04f0a
          20235 => x"81", -- $04f0b
          20236 => x"82", -- $04f0c
          20237 => x"81", -- $04f0d
          20238 => x"81", -- $04f0e
          20239 => x"82", -- $04f0f
          20240 => x"82", -- $04f10
          20241 => x"81", -- $04f11
          20242 => x"82", -- $04f12
          20243 => x"83", -- $04f13
          20244 => x"82", -- $04f14
          20245 => x"82", -- $04f15
          20246 => x"83", -- $04f16
          20247 => x"83", -- $04f17
          20248 => x"83", -- $04f18
          20249 => x"82", -- $04f19
          20250 => x"84", -- $04f1a
          20251 => x"84", -- $04f1b
          20252 => x"82", -- $04f1c
          20253 => x"84", -- $04f1d
          20254 => x"84", -- $04f1e
          20255 => x"84", -- $04f1f
          20256 => x"84", -- $04f20
          20257 => x"84", -- $04f21
          20258 => x"84", -- $04f22
          20259 => x"83", -- $04f23
          20260 => x"83", -- $04f24
          20261 => x"83", -- $04f25
          20262 => x"82", -- $04f26
          20263 => x"81", -- $04f27
          20264 => x"81", -- $04f28
          20265 => x"81", -- $04f29
          20266 => x"80", -- $04f2a
          20267 => x"80", -- $04f2b
          20268 => x"80", -- $04f2c
          20269 => x"80", -- $04f2d
          20270 => x"7f", -- $04f2e
          20271 => x"80", -- $04f2f
          20272 => x"80", -- $04f30
          20273 => x"7f", -- $04f31
          20274 => x"80", -- $04f32
          20275 => x"82", -- $04f33
          20276 => x"82", -- $04f34
          20277 => x"81", -- $04f35
          20278 => x"82", -- $04f36
          20279 => x"83", -- $04f37
          20280 => x"81", -- $04f38
          20281 => x"80", -- $04f39
          20282 => x"81", -- $04f3a
          20283 => x"80", -- $04f3b
          20284 => x"80", -- $04f3c
          20285 => x"7f", -- $04f3d
          20286 => x"80", -- $04f3e
          20287 => x"7f", -- $04f3f
          20288 => x"7e", -- $04f40
          20289 => x"7f", -- $04f41
          20290 => x"7f", -- $04f42
          20291 => x"7f", -- $04f43
          20292 => x"7e", -- $04f44
          20293 => x"7f", -- $04f45
          20294 => x"80", -- $04f46
          20295 => x"80", -- $04f47
          20296 => x"80", -- $04f48
          20297 => x"80", -- $04f49
          20298 => x"81", -- $04f4a
          20299 => x"80", -- $04f4b
          20300 => x"80", -- $04f4c
          20301 => x"81", -- $04f4d
          20302 => x"81", -- $04f4e
          20303 => x"80", -- $04f4f
          20304 => x"80", -- $04f50
          20305 => x"80", -- $04f51
          20306 => x"80", -- $04f52
          20307 => x"80", -- $04f53
          20308 => x"80", -- $04f54
          20309 => x"81", -- $04f55
          20310 => x"80", -- $04f56
          20311 => x"81", -- $04f57
          20312 => x"82", -- $04f58
          20313 => x"82", -- $04f59
          20314 => x"83", -- $04f5a
          20315 => x"84", -- $04f5b
          20316 => x"85", -- $04f5c
          20317 => x"86", -- $04f5d
          20318 => x"87", -- $04f5e
          20319 => x"88", -- $04f5f
          20320 => x"88", -- $04f60
          20321 => x"87", -- $04f61
          20322 => x"89", -- $04f62
          20323 => x"88", -- $04f63
          20324 => x"86", -- $04f64
          20325 => x"88", -- $04f65
          20326 => x"86", -- $04f66
          20327 => x"85", -- $04f67
          20328 => x"83", -- $04f68
          20329 => x"83", -- $04f69
          20330 => x"82", -- $04f6a
          20331 => x"80", -- $04f6b
          20332 => x"7f", -- $04f6c
          20333 => x"7e", -- $04f6d
          20334 => x"7d", -- $04f6e
          20335 => x"7c", -- $04f6f
          20336 => x"7c", -- $04f70
          20337 => x"7b", -- $04f71
          20338 => x"7a", -- $04f72
          20339 => x"7a", -- $04f73
          20340 => x"7b", -- $04f74
          20341 => x"7b", -- $04f75
          20342 => x"7b", -- $04f76
          20343 => x"7c", -- $04f77
          20344 => x"7e", -- $04f78
          20345 => x"7e", -- $04f79
          20346 => x"7f", -- $04f7a
          20347 => x"80", -- $04f7b
          20348 => x"81", -- $04f7c
          20349 => x"82", -- $04f7d
          20350 => x"83", -- $04f7e
          20351 => x"83", -- $04f7f
          20352 => x"83", -- $04f80
          20353 => x"83", -- $04f81
          20354 => x"83", -- $04f82
          20355 => x"82", -- $04f83
          20356 => x"81", -- $04f84
          20357 => x"80", -- $04f85
          20358 => x"7f", -- $04f86
          20359 => x"7e", -- $04f87
          20360 => x"7d", -- $04f88
          20361 => x"7b", -- $04f89
          20362 => x"7c", -- $04f8a
          20363 => x"7c", -- $04f8b
          20364 => x"7b", -- $04f8c
          20365 => x"7c", -- $04f8d
          20366 => x"7d", -- $04f8e
          20367 => x"7d", -- $04f8f
          20368 => x"7d", -- $04f90
          20369 => x"7d", -- $04f91
          20370 => x"7f", -- $04f92
          20371 => x"7f", -- $04f93
          20372 => x"7f", -- $04f94
          20373 => x"80", -- $04f95
          20374 => x"80", -- $04f96
          20375 => x"80", -- $04f97
          20376 => x"80", -- $04f98
          20377 => x"81", -- $04f99
          20378 => x"80", -- $04f9a
          20379 => x"81", -- $04f9b
          20380 => x"82", -- $04f9c
          20381 => x"82", -- $04f9d
          20382 => x"83", -- $04f9e
          20383 => x"83", -- $04f9f
          20384 => x"83", -- $04fa0
          20385 => x"84", -- $04fa1
          20386 => x"83", -- $04fa2
          20387 => x"83", -- $04fa3
          20388 => x"83", -- $04fa4
          20389 => x"82", -- $04fa5
          20390 => x"82", -- $04fa6
          20391 => x"82", -- $04fa7
          20392 => x"81", -- $04fa8
          20393 => x"82", -- $04fa9
          20394 => x"81", -- $04faa
          20395 => x"81", -- $04fab
          20396 => x"82", -- $04fac
          20397 => x"81", -- $04fad
          20398 => x"81", -- $04fae
          20399 => x"81", -- $04faf
          20400 => x"81", -- $04fb0
          20401 => x"81", -- $04fb1
          20402 => x"80", -- $04fb2
          20403 => x"81", -- $04fb3
          20404 => x"80", -- $04fb4
          20405 => x"80", -- $04fb5
          20406 => x"7f", -- $04fb6
          20407 => x"80", -- $04fb7
          20408 => x"7f", -- $04fb8
          20409 => x"7e", -- $04fb9
          20410 => x"80", -- $04fba
          20411 => x"7f", -- $04fbb
          20412 => x"7f", -- $04fbc
          20413 => x"7f", -- $04fbd
          20414 => x"80", -- $04fbe
          20415 => x"80", -- $04fbf
          20416 => x"7f", -- $04fc0
          20417 => x"7f", -- $04fc1
          20418 => x"80", -- $04fc2
          20419 => x"7e", -- $04fc3
          20420 => x"7e", -- $04fc4
          20421 => x"7e", -- $04fc5
          20422 => x"7d", -- $04fc6
          20423 => x"7c", -- $04fc7
          20424 => x"7c", -- $04fc8
          20425 => x"7c", -- $04fc9
          20426 => x"7b", -- $04fca
          20427 => x"7b", -- $04fcb
          20428 => x"7d", -- $04fcc
          20429 => x"7d", -- $04fcd
          20430 => x"7c", -- $04fce
          20431 => x"7e", -- $04fcf
          20432 => x"7e", -- $04fd0
          20433 => x"7e", -- $04fd1
          20434 => x"7f", -- $04fd2
          20435 => x"80", -- $04fd3
          20436 => x"7f", -- $04fd4
          20437 => x"7f", -- $04fd5
          20438 => x"80", -- $04fd6
          20439 => x"7f", -- $04fd7
          20440 => x"7f", -- $04fd8
          20441 => x"7f", -- $04fd9
          20442 => x"80", -- $04fda
          20443 => x"7f", -- $04fdb
          20444 => x"7f", -- $04fdc
          20445 => x"80", -- $04fdd
          20446 => x"7f", -- $04fde
          20447 => x"7f", -- $04fdf
          20448 => x"80", -- $04fe0
          20449 => x"80", -- $04fe1
          20450 => x"80", -- $04fe2
          20451 => x"80", -- $04fe3
          20452 => x"81", -- $04fe4
          20453 => x"81", -- $04fe5
          20454 => x"81", -- $04fe6
          20455 => x"83", -- $04fe7
          20456 => x"83", -- $04fe8
          20457 => x"83", -- $04fe9
          20458 => x"84", -- $04fea
          20459 => x"85", -- $04feb
          20460 => x"85", -- $04fec
          20461 => x"85", -- $04fed
          20462 => x"85", -- $04fee
          20463 => x"84", -- $04fef
          20464 => x"85", -- $04ff0
          20465 => x"83", -- $04ff1
          20466 => x"83", -- $04ff2
          20467 => x"84", -- $04ff3
          20468 => x"81", -- $04ff4
          20469 => x"81", -- $04ff5
          20470 => x"81", -- $04ff6
          20471 => x"80", -- $04ff7
          20472 => x"80", -- $04ff8
          20473 => x"7f", -- $04ff9
          20474 => x"7f", -- $04ffa
          20475 => x"7e", -- $04ffb
          20476 => x"7d", -- $04ffc
          20477 => x"7c", -- $04ffd
          20478 => x"7c", -- $04ffe
          20479 => x"7b", -- $04fff
          20480 => x"7a", -- $05000
          20481 => x"7a", -- $05001
          20482 => x"7a", -- $05002
          20483 => x"7a", -- $05003
          20484 => x"7a", -- $05004
          20485 => x"7b", -- $05005
          20486 => x"7b", -- $05006
          20487 => x"7b", -- $05007
          20488 => x"7d", -- $05008
          20489 => x"7e", -- $05009
          20490 => x"7f", -- $0500a
          20491 => x"80", -- $0500b
          20492 => x"80", -- $0500c
          20493 => x"80", -- $0500d
          20494 => x"80", -- $0500e
          20495 => x"80", -- $0500f
          20496 => x"80", -- $05010
          20497 => x"7f", -- $05011
          20498 => x"7e", -- $05012
          20499 => x"7e", -- $05013
          20500 => x"7d", -- $05014
          20501 => x"7c", -- $05015
          20502 => x"7c", -- $05016
          20503 => x"7c", -- $05017
          20504 => x"7b", -- $05018
          20505 => x"7b", -- $05019
          20506 => x"7c", -- $0501a
          20507 => x"7d", -- $0501b
          20508 => x"7d", -- $0501c
          20509 => x"7e", -- $0501d
          20510 => x"7f", -- $0501e
          20511 => x"7f", -- $0501f
          20512 => x"80", -- $05020
          20513 => x"80", -- $05021
          20514 => x"80", -- $05022
          20515 => x"80", -- $05023
          20516 => x"81", -- $05024
          20517 => x"82", -- $05025
          20518 => x"82", -- $05026
          20519 => x"82", -- $05027
          20520 => x"82", -- $05028
          20521 => x"83", -- $05029
          20522 => x"82", -- $0502a
          20523 => x"83", -- $0502b
          20524 => x"83", -- $0502c
          20525 => x"83", -- $0502d
          20526 => x"84", -- $0502e
          20527 => x"83", -- $0502f
          20528 => x"83", -- $05030
          20529 => x"84", -- $05031
          20530 => x"83", -- $05032
          20531 => x"83", -- $05033
          20532 => x"84", -- $05034
          20533 => x"84", -- $05035
          20534 => x"84", -- $05036
          20535 => x"84", -- $05037
          20536 => x"83", -- $05038
          20537 => x"83", -- $05039
          20538 => x"82", -- $0503a
          20539 => x"80", -- $0503b
          20540 => x"80", -- $0503c
          20541 => x"7f", -- $0503d
          20542 => x"7f", -- $0503e
          20543 => x"7e", -- $0503f
          20544 => x"7c", -- $05040
          20545 => x"7b", -- $05041
          20546 => x"7b", -- $05042
          20547 => x"7a", -- $05043
          20548 => x"7a", -- $05044
          20549 => x"7a", -- $05045
          20550 => x"7a", -- $05046
          20551 => x"7a", -- $05047
          20552 => x"7b", -- $05048
          20553 => x"7b", -- $05049
          20554 => x"7b", -- $0504a
          20555 => x"7c", -- $0504b
          20556 => x"7c", -- $0504c
          20557 => x"7d", -- $0504d
          20558 => x"7d", -- $0504e
          20559 => x"7e", -- $0504f
          20560 => x"7e", -- $05050
          20561 => x"7e", -- $05051
          20562 => x"7f", -- $05052
          20563 => x"7f", -- $05053
          20564 => x"7f", -- $05054
          20565 => x"7e", -- $05055
          20566 => x"7e", -- $05056
          20567 => x"7e", -- $05057
          20568 => x"7d", -- $05058
          20569 => x"7c", -- $05059
          20570 => x"7c", -- $0505a
          20571 => x"7c", -- $0505b
          20572 => x"7b", -- $0505c
          20573 => x"7c", -- $0505d
          20574 => x"7c", -- $0505e
          20575 => x"7c", -- $0505f
          20576 => x"7d", -- $05060
          20577 => x"7e", -- $05061
          20578 => x"7f", -- $05062
          20579 => x"80", -- $05063
          20580 => x"80", -- $05064
          20581 => x"80", -- $05065
          20582 => x"81", -- $05066
          20583 => x"81", -- $05067
          20584 => x"82", -- $05068
          20585 => x"83", -- $05069
          20586 => x"82", -- $0506a
          20587 => x"83", -- $0506b
          20588 => x"83", -- $0506c
          20589 => x"82", -- $0506d
          20590 => x"82", -- $0506e
          20591 => x"82", -- $0506f
          20592 => x"81", -- $05070
          20593 => x"82", -- $05071
          20594 => x"83", -- $05072
          20595 => x"83", -- $05073
          20596 => x"84", -- $05074
          20597 => x"85", -- $05075
          20598 => x"85", -- $05076
          20599 => x"86", -- $05077
          20600 => x"85", -- $05078
          20601 => x"85", -- $05079
          20602 => x"85", -- $0507a
          20603 => x"83", -- $0507b
          20604 => x"83", -- $0507c
          20605 => x"82", -- $0507d
          20606 => x"80", -- $0507e
          20607 => x"80", -- $0507f
          20608 => x"7f", -- $05080
          20609 => x"7e", -- $05081
          20610 => x"7c", -- $05082
          20611 => x"7c", -- $05083
          20612 => x"7b", -- $05084
          20613 => x"7a", -- $05085
          20614 => x"79", -- $05086
          20615 => x"78", -- $05087
          20616 => x"78", -- $05088
          20617 => x"77", -- $05089
          20618 => x"77", -- $0508a
          20619 => x"78", -- $0508b
          20620 => x"78", -- $0508c
          20621 => x"79", -- $0508d
          20622 => x"7a", -- $0508e
          20623 => x"7a", -- $0508f
          20624 => x"7b", -- $05090
          20625 => x"7c", -- $05091
          20626 => x"7d", -- $05092
          20627 => x"7e", -- $05093
          20628 => x"7e", -- $05094
          20629 => x"7f", -- $05095
          20630 => x"7e", -- $05096
          20631 => x"7e", -- $05097
          20632 => x"7e", -- $05098
          20633 => x"7d", -- $05099
          20634 => x"7c", -- $0509a
          20635 => x"7b", -- $0509b
          20636 => x"7a", -- $0509c
          20637 => x"7a", -- $0509d
          20638 => x"7a", -- $0509e
          20639 => x"7a", -- $0509f
          20640 => x"7a", -- $050a0
          20641 => x"7b", -- $050a1
          20642 => x"7b", -- $050a2
          20643 => x"7c", -- $050a3
          20644 => x"7e", -- $050a4
          20645 => x"7e", -- $050a5
          20646 => x"7f", -- $050a6
          20647 => x"80", -- $050a7
          20648 => x"80", -- $050a8
          20649 => x"80", -- $050a9
          20650 => x"81", -- $050aa
          20651 => x"81", -- $050ab
          20652 => x"81", -- $050ac
          20653 => x"81", -- $050ad
          20654 => x"81", -- $050ae
          20655 => x"82", -- $050af
          20656 => x"82", -- $050b0
          20657 => x"82", -- $050b1
          20658 => x"83", -- $050b2
          20659 => x"83", -- $050b3
          20660 => x"84", -- $050b4
          20661 => x"85", -- $050b5
          20662 => x"86", -- $050b6
          20663 => x"86", -- $050b7
          20664 => x"86", -- $050b8
          20665 => x"87", -- $050b9
          20666 => x"86", -- $050ba
          20667 => x"86", -- $050bb
          20668 => x"86", -- $050bc
          20669 => x"85", -- $050bd
          20670 => x"84", -- $050be
          20671 => x"83", -- $050bf
          20672 => x"83", -- $050c0
          20673 => x"82", -- $050c1
          20674 => x"80", -- $050c2
          20675 => x"80", -- $050c3
          20676 => x"7e", -- $050c4
          20677 => x"7c", -- $050c5
          20678 => x"7b", -- $050c6
          20679 => x"7a", -- $050c7
          20680 => x"79", -- $050c8
          20681 => x"78", -- $050c9
          20682 => x"78", -- $050ca
          20683 => x"78", -- $050cb
          20684 => x"78", -- $050cc
          20685 => x"78", -- $050cd
          20686 => x"79", -- $050ce
          20687 => x"7a", -- $050cf
          20688 => x"7b", -- $050d0
          20689 => x"7c", -- $050d1
          20690 => x"7d", -- $050d2
          20691 => x"7e", -- $050d3
          20692 => x"7f", -- $050d4
          20693 => x"80", -- $050d5
          20694 => x"80", -- $050d6
          20695 => x"80", -- $050d7
          20696 => x"80", -- $050d8
          20697 => x"7f", -- $050d9
          20698 => x"7f", -- $050da
          20699 => x"7e", -- $050db
          20700 => x"7e", -- $050dc
          20701 => x"7d", -- $050dd
          20702 => x"7d", -- $050de
          20703 => x"7d", -- $050df
          20704 => x"7d", -- $050e0
          20705 => x"7d", -- $050e1
          20706 => x"7d", -- $050e2
          20707 => x"7d", -- $050e3
          20708 => x"7e", -- $050e4
          20709 => x"7f", -- $050e5
          20710 => x"80", -- $050e6
          20711 => x"80", -- $050e7
          20712 => x"80", -- $050e8
          20713 => x"81", -- $050e9
          20714 => x"81", -- $050ea
          20715 => x"82", -- $050eb
          20716 => x"83", -- $050ec
          20717 => x"83", -- $050ed
          20718 => x"84", -- $050ee
          20719 => x"84", -- $050ef
          20720 => x"84", -- $050f0
          20721 => x"84", -- $050f1
          20722 => x"84", -- $050f2
          20723 => x"84", -- $050f3
          20724 => x"84", -- $050f4
          20725 => x"85", -- $050f5
          20726 => x"85", -- $050f6
          20727 => x"86", -- $050f7
          20728 => x"87", -- $050f8
          20729 => x"86", -- $050f9
          20730 => x"88", -- $050fa
          20731 => x"88", -- $050fb
          20732 => x"88", -- $050fc
          20733 => x"88", -- $050fd
          20734 => x"87", -- $050fe
          20735 => x"87", -- $050ff
          20736 => x"86", -- $05100
          20737 => x"85", -- $05101
          20738 => x"85", -- $05102
          20739 => x"83", -- $05103
          20740 => x"82", -- $05104
          20741 => x"81", -- $05105
          20742 => x"80", -- $05106
          20743 => x"7f", -- $05107
          20744 => x"7d", -- $05108
          20745 => x"7d", -- $05109
          20746 => x"7c", -- $0510a
          20747 => x"7b", -- $0510b
          20748 => x"7b", -- $0510c
          20749 => x"7a", -- $0510d
          20750 => x"7a", -- $0510e
          20751 => x"7a", -- $0510f
          20752 => x"7b", -- $05110
          20753 => x"7b", -- $05111
          20754 => x"7c", -- $05112
          20755 => x"7c", -- $05113
          20756 => x"7d", -- $05114
          20757 => x"7d", -- $05115
          20758 => x"7d", -- $05116
          20759 => x"7d", -- $05117
          20760 => x"7e", -- $05118
          20761 => x"7e", -- $05119
          20762 => x"7e", -- $0511a
          20763 => x"7e", -- $0511b
          20764 => x"7e", -- $0511c
          20765 => x"7e", -- $0511d
          20766 => x"7d", -- $0511e
          20767 => x"7d", -- $0511f
          20768 => x"7d", -- $05120
          20769 => x"7d", -- $05121
          20770 => x"7d", -- $05122
          20771 => x"7e", -- $05123
          20772 => x"7e", -- $05124
          20773 => x"7e", -- $05125
          20774 => x"7e", -- $05126
          20775 => x"7f", -- $05127
          20776 => x"80", -- $05128
          20777 => x"80", -- $05129
          20778 => x"81", -- $0512a
          20779 => x"82", -- $0512b
          20780 => x"83", -- $0512c
          20781 => x"84", -- $0512d
          20782 => x"85", -- $0512e
          20783 => x"85", -- $0512f
          20784 => x"86", -- $05130
          20785 => x"86", -- $05131
          20786 => x"86", -- $05132
          20787 => x"86", -- $05133
          20788 => x"87", -- $05134
          20789 => x"86", -- $05135
          20790 => x"86", -- $05136
          20791 => x"86", -- $05137
          20792 => x"87", -- $05138
          20793 => x"87", -- $05139
          20794 => x"87", -- $0513a
          20795 => x"88", -- $0513b
          20796 => x"87", -- $0513c
          20797 => x"88", -- $0513d
          20798 => x"87", -- $0513e
          20799 => x"86", -- $0513f
          20800 => x"86", -- $05140
          20801 => x"85", -- $05141
          20802 => x"84", -- $05142
          20803 => x"83", -- $05143
          20804 => x"83", -- $05144
          20805 => x"81", -- $05145
          20806 => x"80", -- $05146
          20807 => x"80", -- $05147
          20808 => x"7f", -- $05148
          20809 => x"7e", -- $05149
          20810 => x"7c", -- $0514a
          20811 => x"7c", -- $0514b
          20812 => x"7b", -- $0514c
          20813 => x"7a", -- $0514d
          20814 => x"7a", -- $0514e
          20815 => x"7a", -- $0514f
          20816 => x"7a", -- $05150
          20817 => x"7a", -- $05151
          20818 => x"7b", -- $05152
          20819 => x"7c", -- $05153
          20820 => x"7b", -- $05154
          20821 => x"7d", -- $05155
          20822 => x"7d", -- $05156
          20823 => x"7d", -- $05157
          20824 => x"7e", -- $05158
          20825 => x"7e", -- $05159
          20826 => x"7e", -- $0515a
          20827 => x"7e", -- $0515b
          20828 => x"7e", -- $0515c
          20829 => x"7e", -- $0515d
          20830 => x"7e", -- $0515e
          20831 => x"7e", -- $0515f
          20832 => x"7d", -- $05160
          20833 => x"7d", -- $05161
          20834 => x"7c", -- $05162
          20835 => x"7d", -- $05163
          20836 => x"7d", -- $05164
          20837 => x"7d", -- $05165
          20838 => x"7d", -- $05166
          20839 => x"7e", -- $05167
          20840 => x"7e", -- $05168
          20841 => x"7f", -- $05169
          20842 => x"80", -- $0516a
          20843 => x"80", -- $0516b
          20844 => x"81", -- $0516c
          20845 => x"83", -- $0516d
          20846 => x"84", -- $0516e
          20847 => x"85", -- $0516f
          20848 => x"85", -- $05170
          20849 => x"86", -- $05171
          20850 => x"86", -- $05172
          20851 => x"87", -- $05173
          20852 => x"87", -- $05174
          20853 => x"87", -- $05175
          20854 => x"87", -- $05176
          20855 => x"87", -- $05177
          20856 => x"88", -- $05178
          20857 => x"87", -- $05179
          20858 => x"88", -- $0517a
          20859 => x"88", -- $0517b
          20860 => x"88", -- $0517c
          20861 => x"88", -- $0517d
          20862 => x"87", -- $0517e
          20863 => x"87", -- $0517f
          20864 => x"86", -- $05180
          20865 => x"86", -- $05181
          20866 => x"86", -- $05182
          20867 => x"85", -- $05183
          20868 => x"85", -- $05184
          20869 => x"84", -- $05185
          20870 => x"83", -- $05186
          20871 => x"82", -- $05187
          20872 => x"81", -- $05188
          20873 => x"80", -- $05189
          20874 => x"80", -- $0518a
          20875 => x"7f", -- $0518b
          20876 => x"7e", -- $0518c
          20877 => x"7d", -- $0518d
          20878 => x"7c", -- $0518e
          20879 => x"7c", -- $0518f
          20880 => x"7c", -- $05190
          20881 => x"7c", -- $05191
          20882 => x"7c", -- $05192
          20883 => x"7c", -- $05193
          20884 => x"7c", -- $05194
          20885 => x"7d", -- $05195
          20886 => x"7e", -- $05196
          20887 => x"7f", -- $05197
          20888 => x"7f", -- $05198
          20889 => x"80", -- $05199
          20890 => x"80", -- $0519a
          20891 => x"80", -- $0519b
          20892 => x"80", -- $0519c
          20893 => x"80", -- $0519d
          20894 => x"80", -- $0519e
          20895 => x"80", -- $0519f
          20896 => x"7f", -- $051a0
          20897 => x"7f", -- $051a1
          20898 => x"7f", -- $051a2
          20899 => x"7e", -- $051a3
          20900 => x"7f", -- $051a4
          20901 => x"7f", -- $051a5
          20902 => x"7f", -- $051a6
          20903 => x"80", -- $051a7
          20904 => x"80", -- $051a8
          20905 => x"80", -- $051a9
          20906 => x"81", -- $051aa
          20907 => x"82", -- $051ab
          20908 => x"82", -- $051ac
          20909 => x"84", -- $051ad
          20910 => x"84", -- $051ae
          20911 => x"85", -- $051af
          20912 => x"86", -- $051b0
          20913 => x"86", -- $051b1
          20914 => x"86", -- $051b2
          20915 => x"86", -- $051b3
          20916 => x"87", -- $051b4
          20917 => x"87", -- $051b5
          20918 => x"87", -- $051b6
          20919 => x"87", -- $051b7
          20920 => x"87", -- $051b8
          20921 => x"87", -- $051b9
          20922 => x"87", -- $051ba
          20923 => x"87", -- $051bb
          20924 => x"87", -- $051bc
          20925 => x"87", -- $051bd
          20926 => x"87", -- $051be
          20927 => x"87", -- $051bf
          20928 => x"87", -- $051c0
          20929 => x"87", -- $051c1
          20930 => x"86", -- $051c2
          20931 => x"86", -- $051c3
          20932 => x"86", -- $051c4
          20933 => x"85", -- $051c5
          20934 => x"84", -- $051c6
          20935 => x"83", -- $051c7
          20936 => x"83", -- $051c8
          20937 => x"81", -- $051c9
          20938 => x"80", -- $051ca
          20939 => x"80", -- $051cb
          20940 => x"7f", -- $051cc
          20941 => x"7e", -- $051cd
          20942 => x"7d", -- $051ce
          20943 => x"7d", -- $051cf
          20944 => x"7c", -- $051d0
          20945 => x"7c", -- $051d1
          20946 => x"7d", -- $051d2
          20947 => x"7d", -- $051d3
          20948 => x"7c", -- $051d4
          20949 => x"7d", -- $051d5
          20950 => x"7d", -- $051d6
          20951 => x"7d", -- $051d7
          20952 => x"7e", -- $051d8
          20953 => x"7e", -- $051d9
          20954 => x"7e", -- $051da
          20955 => x"7e", -- $051db
          20956 => x"7e", -- $051dc
          20957 => x"7f", -- $051dd
          20958 => x"7f", -- $051de
          20959 => x"7f", -- $051df
          20960 => x"7e", -- $051e0
          20961 => x"7e", -- $051e1
          20962 => x"7e", -- $051e2
          20963 => x"7e", -- $051e3
          20964 => x"7e", -- $051e4
          20965 => x"7e", -- $051e5
          20966 => x"7e", -- $051e6
          20967 => x"7f", -- $051e7
          20968 => x"80", -- $051e8
          20969 => x"80", -- $051e9
          20970 => x"80", -- $051ea
          20971 => x"80", -- $051eb
          20972 => x"81", -- $051ec
          20973 => x"81", -- $051ed
          20974 => x"83", -- $051ee
          20975 => x"84", -- $051ef
          20976 => x"84", -- $051f0
          20977 => x"86", -- $051f1
          20978 => x"87", -- $051f2
          20979 => x"86", -- $051f3
          20980 => x"87", -- $051f4
          20981 => x"87", -- $051f5
          20982 => x"87", -- $051f6
          20983 => x"88", -- $051f7
          20984 => x"87", -- $051f8
          20985 => x"87", -- $051f9
          20986 => x"87", -- $051fa
          20987 => x"86", -- $051fb
          20988 => x"87", -- $051fc
          20989 => x"86", -- $051fd
          20990 => x"86", -- $051fe
          20991 => x"86", -- $051ff
          20992 => x"86", -- $05200
          20993 => x"85", -- $05201
          20994 => x"84", -- $05202
          20995 => x"84", -- $05203
          20996 => x"83", -- $05204
          20997 => x"83", -- $05205
          20998 => x"82", -- $05206
          20999 => x"82", -- $05207
          21000 => x"81", -- $05208
          21001 => x"81", -- $05209
          21002 => x"80", -- $0520a
          21003 => x"80", -- $0520b
          21004 => x"80", -- $0520c
          21005 => x"80", -- $0520d
          21006 => x"80", -- $0520e
          21007 => x"80", -- $0520f
          21008 => x"80", -- $05210
          21009 => x"80", -- $05211
          21010 => x"80", -- $05212
          21011 => x"80", -- $05213
          21012 => x"80", -- $05214
          21013 => x"80", -- $05215
          21014 => x"80", -- $05216
          21015 => x"80", -- $05217
          21016 => x"80", -- $05218
          21017 => x"80", -- $05219
          21018 => x"7f", -- $0521a
          21019 => x"7f", -- $0521b
          21020 => x"7e", -- $0521c
          21021 => x"7e", -- $0521d
          21022 => x"7d", -- $0521e
          21023 => x"7d", -- $0521f
          21024 => x"7c", -- $05220
          21025 => x"7c", -- $05221
          21026 => x"7c", -- $05222
          21027 => x"7c", -- $05223
          21028 => x"7c", -- $05224
          21029 => x"7c", -- $05225
          21030 => x"7c", -- $05226
          21031 => x"7d", -- $05227
          21032 => x"7e", -- $05228
          21033 => x"7e", -- $05229
          21034 => x"7f", -- $0522a
          21035 => x"80", -- $0522b
          21036 => x"80", -- $0522c
          21037 => x"80", -- $0522d
          21038 => x"81", -- $0522e
          21039 => x"82", -- $0522f
          21040 => x"83", -- $05230
          21041 => x"83", -- $05231
          21042 => x"84", -- $05232
          21043 => x"85", -- $05233
          21044 => x"85", -- $05234
          21045 => x"85", -- $05235
          21046 => x"86", -- $05236
          21047 => x"86", -- $05237
          21048 => x"87", -- $05238
          21049 => x"86", -- $05239
          21050 => x"86", -- $0523a
          21051 => x"86", -- $0523b
          21052 => x"85", -- $0523c
          21053 => x"85", -- $0523d
          21054 => x"84", -- $0523e
          21055 => x"84", -- $0523f
          21056 => x"83", -- $05240
          21057 => x"83", -- $05241
          21058 => x"82", -- $05242
          21059 => x"81", -- $05243
          21060 => x"80", -- $05244
          21061 => x"80", -- $05245
          21062 => x"80", -- $05246
          21063 => x"80", -- $05247
          21064 => x"7f", -- $05248
          21065 => x"7f", -- $05249
          21066 => x"7f", -- $0524a
          21067 => x"7e", -- $0524b
          21068 => x"7e", -- $0524c
          21069 => x"7e", -- $0524d
          21070 => x"7e", -- $0524e
          21071 => x"7e", -- $0524f
          21072 => x"7e", -- $05250
          21073 => x"7e", -- $05251
          21074 => x"7e", -- $05252
          21075 => x"7e", -- $05253
          21076 => x"7e", -- $05254
          21077 => x"7e", -- $05255
          21078 => x"7e", -- $05256
          21079 => x"7e", -- $05257
          21080 => x"7e", -- $05258
          21081 => x"7e", -- $05259
          21082 => x"7e", -- $0525a
          21083 => x"7d", -- $0525b
          21084 => x"7d", -- $0525c
          21085 => x"7d", -- $0525d
          21086 => x"7d", -- $0525e
          21087 => x"7c", -- $0525f
          21088 => x"7c", -- $05260
          21089 => x"7c", -- $05261
          21090 => x"7c", -- $05262
          21091 => x"7c", -- $05263
          21092 => x"7c", -- $05264
          21093 => x"7c", -- $05265
          21094 => x"7d", -- $05266
          21095 => x"7d", -- $05267
          21096 => x"7e", -- $05268
          21097 => x"7e", -- $05269
          21098 => x"7e", -- $0526a
          21099 => x"7f", -- $0526b
          21100 => x"7f", -- $0526c
          21101 => x"80", -- $0526d
          21102 => x"80", -- $0526e
          21103 => x"80", -- $0526f
          21104 => x"81", -- $05270
          21105 => x"81", -- $05271
          21106 => x"81", -- $05272
          21107 => x"82", -- $05273
          21108 => x"82", -- $05274
          21109 => x"83", -- $05275
          21110 => x"83", -- $05276
          21111 => x"82", -- $05277
          21112 => x"83", -- $05278
          21113 => x"83", -- $05279
          21114 => x"82", -- $0527a
          21115 => x"82", -- $0527b
          21116 => x"83", -- $0527c
          21117 => x"83", -- $0527d
          21118 => x"82", -- $0527e
          21119 => x"82", -- $0527f
          21120 => x"81", -- $05280
          21121 => x"81", -- $05281
          21122 => x"80", -- $05282
          21123 => x"80", -- $05283
          21124 => x"80", -- $05284
          21125 => x"80", -- $05285
          21126 => x"80", -- $05286
          21127 => x"80", -- $05287
          21128 => x"80", -- $05288
          21129 => x"80", -- $05289
          21130 => x"80", -- $0528a
          21131 => x"7f", -- $0528b
          21132 => x"7f", -- $0528c
          21133 => x"7f", -- $0528d
          21134 => x"7e", -- $0528e
          21135 => x"7f", -- $0528f
          21136 => x"7f", -- $05290
          21137 => x"7e", -- $05291
          21138 => x"7e", -- $05292
          21139 => x"7e", -- $05293
          21140 => x"7d", -- $05294
          21141 => x"7d", -- $05295
          21142 => x"7c", -- $05296
          21143 => x"7c", -- $05297
          21144 => x"7c", -- $05298
          21145 => x"7c", -- $05299
          21146 => x"7b", -- $0529a
          21147 => x"7b", -- $0529b
          21148 => x"7b", -- $0529c
          21149 => x"7b", -- $0529d
          21150 => x"7b", -- $0529e
          21151 => x"7b", -- $0529f
          21152 => x"7b", -- $052a0
          21153 => x"7c", -- $052a1
          21154 => x"7c", -- $052a2
          21155 => x"7c", -- $052a3
          21156 => x"7c", -- $052a4
          21157 => x"7d", -- $052a5
          21158 => x"7d", -- $052a6
          21159 => x"7e", -- $052a7
          21160 => x"7f", -- $052a8
          21161 => x"7f", -- $052a9
          21162 => x"7f", -- $052aa
          21163 => x"80", -- $052ab
          21164 => x"80", -- $052ac
          21165 => x"81", -- $052ad
          21166 => x"81", -- $052ae
          21167 => x"81", -- $052af
          21168 => x"82", -- $052b0
          21169 => x"82", -- $052b1
          21170 => x"82", -- $052b2
          21171 => x"82", -- $052b3
          21172 => x"83", -- $052b4
          21173 => x"84", -- $052b5
          21174 => x"83", -- $052b6
          21175 => x"83", -- $052b7
          21176 => x"83", -- $052b8
          21177 => x"83", -- $052b9
          21178 => x"82", -- $052ba
          21179 => x"82", -- $052bb
          21180 => x"82", -- $052bc
          21181 => x"81", -- $052bd
          21182 => x"80", -- $052be
          21183 => x"80", -- $052bf
          21184 => x"80", -- $052c0
          21185 => x"80", -- $052c1
          21186 => x"80", -- $052c2
          21187 => x"80", -- $052c3
          21188 => x"7f", -- $052c4
          21189 => x"7f", -- $052c5
          21190 => x"7f", -- $052c6
          21191 => x"7e", -- $052c7
          21192 => x"7e", -- $052c8
          21193 => x"7f", -- $052c9
          21194 => x"7f", -- $052ca
          21195 => x"7f", -- $052cb
          21196 => x"7f", -- $052cc
          21197 => x"7f", -- $052cd
          21198 => x"7f", -- $052ce
          21199 => x"7f", -- $052cf
          21200 => x"7e", -- $052d0
          21201 => x"7e", -- $052d1
          21202 => x"7e", -- $052d2
          21203 => x"7d", -- $052d3
          21204 => x"7d", -- $052d4
          21205 => x"7e", -- $052d5
          21206 => x"7e", -- $052d6
          21207 => x"7e", -- $052d7
          21208 => x"7e", -- $052d8
          21209 => x"7e", -- $052d9
          21210 => x"7e", -- $052da
          21211 => x"7e", -- $052db
          21212 => x"7d", -- $052dc
          21213 => x"7d", -- $052dd
          21214 => x"7d", -- $052de
          21215 => x"7d", -- $052df
          21216 => x"7d", -- $052e0
          21217 => x"7d", -- $052e1
          21218 => x"7d", -- $052e2
          21219 => x"7d", -- $052e3
          21220 => x"7d", -- $052e4
          21221 => x"7d", -- $052e5
          21222 => x"7d", -- $052e6
          21223 => x"7d", -- $052e7
          21224 => x"7d", -- $052e8
          21225 => x"7d", -- $052e9
          21226 => x"7e", -- $052ea
          21227 => x"7e", -- $052eb
          21228 => x"7f", -- $052ec
          21229 => x"7f", -- $052ed
          21230 => x"7f", -- $052ee
          21231 => x"7f", -- $052ef
          21232 => x"7f", -- $052f0
          21233 => x"7f", -- $052f1
          21234 => x"7f", -- $052f2
          21235 => x"7f", -- $052f3
          21236 => x"80", -- $052f4
          21237 => x"80", -- $052f5
          21238 => x"80", -- $052f6
          21239 => x"81", -- $052f7
          21240 => x"81", -- $052f8
          21241 => x"81", -- $052f9
          21242 => x"81", -- $052fa
          21243 => x"80", -- $052fb
          21244 => x"80", -- $052fc
          21245 => x"80", -- $052fd
          21246 => x"80", -- $052fe
          21247 => x"80", -- $052ff
          21248 => x"80", -- $05300
          21249 => x"80", -- $05301
          21250 => x"80", -- $05302
          21251 => x"7f", -- $05303
          21252 => x"7f", -- $05304
          21253 => x"7f", -- $05305
          21254 => x"7e", -- $05306
          21255 => x"7e", -- $05307
          21256 => x"7e", -- $05308
          21257 => x"7d", -- $05309
          21258 => x"7d", -- $0530a
          21259 => x"7d", -- $0530b
          21260 => x"7d", -- $0530c
          21261 => x"7d", -- $0530d
          21262 => x"7c", -- $0530e
          21263 => x"7c", -- $0530f
          21264 => x"7c", -- $05310
          21265 => x"7c", -- $05311
          21266 => x"7c", -- $05312
          21267 => x"7d", -- $05313
          21268 => x"7d", -- $05314
          21269 => x"7d", -- $05315
          21270 => x"7d", -- $05316
          21271 => x"7d", -- $05317
          21272 => x"7c", -- $05318
          21273 => x"7c", -- $05319
          21274 => x"7c", -- $0531a
          21275 => x"7d", -- $0531b
          21276 => x"7e", -- $0531c
          21277 => x"7e", -- $0531d
          21278 => x"7e", -- $0531e
          21279 => x"7e", -- $0531f
          21280 => x"7e", -- $05320
          21281 => x"7e", -- $05321
          21282 => x"7e", -- $05322
          21283 => x"7e", -- $05323
          21284 => x"7e", -- $05324
          21285 => x"7e", -- $05325
          21286 => x"7e", -- $05326
          21287 => x"7f", -- $05327
          21288 => x"7f", -- $05328
          21289 => x"7f", -- $05329
          21290 => x"7f", -- $0532a
          21291 => x"7f", -- $0532b
          21292 => x"7f", -- $0532c
          21293 => x"80", -- $0532d
          21294 => x"80", -- $0532e
          21295 => x"80", -- $0532f
          21296 => x"80", -- $05330
          21297 => x"80", -- $05331
          21298 => x"80", -- $05332
          21299 => x"80", -- $05333
          21300 => x"80", -- $05334
          21301 => x"80", -- $05335
          21302 => x"80", -- $05336
          21303 => x"80", -- $05337
          21304 => x"80", -- $05338
          21305 => x"80", -- $05339
          21306 => x"80", -- $0533a
          21307 => x"80", -- $0533b
          21308 => x"80", -- $0533c
          21309 => x"80", -- $0533d
          21310 => x"80", -- $0533e
          21311 => x"80", -- $0533f
          21312 => x"80", -- $05340
          21313 => x"80", -- $05341
          21314 => x"80", -- $05342
          21315 => x"80", -- $05343
          21316 => x"80", -- $05344
          21317 => x"80", -- $05345
          21318 => x"80", -- $05346
          21319 => x"80", -- $05347
          21320 => x"7f", -- $05348
          21321 => x"7f", -- $05349
          21322 => x"7f", -- $0534a
          21323 => x"7f", -- $0534b
          21324 => x"7f", -- $0534c
          21325 => x"7e", -- $0534d
          21326 => x"7e", -- $0534e
          21327 => x"7e", -- $0534f
          21328 => x"7e", -- $05350
          21329 => x"7e", -- $05351
          21330 => x"7e", -- $05352
          21331 => x"7e", -- $05353
          21332 => x"7e", -- $05354
          21333 => x"7f", -- $05355
          21334 => x"7e", -- $05356
          21335 => x"7e", -- $05357
          21336 => x"7e", -- $05358
          21337 => x"7d", -- $05359
          21338 => x"7d", -- $0535a
          21339 => x"7d", -- $0535b
          21340 => x"7c", -- $0535c
          21341 => x"7d", -- $0535d
          21342 => x"7d", -- $0535e
          21343 => x"7d", -- $0535f
          21344 => x"7e", -- $05360
          21345 => x"7e", -- $05361
          21346 => x"7e", -- $05362
          21347 => x"7e", -- $05363
          21348 => x"7f", -- $05364
          21349 => x"7f", -- $05365
          21350 => x"7f", -- $05366
          21351 => x"7f", -- $05367
          21352 => x"80", -- $05368
          21353 => x"80", -- $05369
          21354 => x"80", -- $0536a
          21355 => x"80", -- $0536b
          21356 => x"80", -- $0536c
          21357 => x"80", -- $0536d
          21358 => x"80", -- $0536e
          21359 => x"80", -- $0536f
          21360 => x"80", -- $05370
          21361 => x"80", -- $05371
          21362 => x"80", -- $05372
          21363 => x"81", -- $05373
          21364 => x"81", -- $05374
          21365 => x"81", -- $05375
          21366 => x"81", -- $05376
          21367 => x"80", -- $05377
          21368 => x"80", -- $05378
          21369 => x"80", -- $05379
          21370 => x"80", -- $0537a
          21371 => x"80", -- $0537b
          21372 => x"80", -- $0537c
          21373 => x"80", -- $0537d
          21374 => x"80", -- $0537e
          21375 => x"80", -- $0537f
          21376 => x"7f", -- $05380
          21377 => x"7f", -- $05381
          21378 => x"7f", -- $05382
          21379 => x"7f", -- $05383
          21380 => x"7f", -- $05384
          21381 => x"7f", -- $05385
          21382 => x"7f", -- $05386
          21383 => x"7f", -- $05387
          21384 => x"80", -- $05388
          21385 => x"7f", -- $05389
          21386 => x"7f", -- $0538a
          21387 => x"7f", -- $0538b
          21388 => x"7e", -- $0538c
          21389 => x"7e", -- $0538d
          21390 => x"7e", -- $0538e
          21391 => x"7e", -- $0538f
          21392 => x"7e", -- $05390
          21393 => x"7f", -- $05391
          21394 => x"7f", -- $05392
          21395 => x"7f", -- $05393
          21396 => x"7f", -- $05394
          21397 => x"7f", -- $05395
          21398 => x"7f", -- $05396
          21399 => x"7f", -- $05397
          21400 => x"7f", -- $05398
          21401 => x"80", -- $05399
          21402 => x"80", -- $0539a
          21403 => x"7f", -- $0539b
          21404 => x"80", -- $0539c
          21405 => x"80", -- $0539d
          21406 => x"80", -- $0539e
          21407 => x"80", -- $0539f
          21408 => x"80", -- $053a0
          21409 => x"80", -- $053a1
          21410 => x"80", -- $053a2
          21411 => x"80", -- $053a3
          21412 => x"80", -- $053a4
          21413 => x"80", -- $053a5
          21414 => x"80", -- $053a6
          21415 => x"80", -- $053a7
          21416 => x"80", -- $053a8
          21417 => x"80", -- $053a9
          21418 => x"80", -- $053aa
          21419 => x"80", -- $053ab
          21420 => x"80", -- $053ac
          21421 => x"80", -- $053ad
          21422 => x"80", -- $053ae
          21423 => x"80", -- $053af
          21424 => x"80", -- $053b0
          21425 => x"80", -- $053b1
          21426 => x"80", -- $053b2
          21427 => x"80", -- $053b3
          21428 => x"80", -- $053b4
          21429 => x"80", -- $053b5
          21430 => x"81", -- $053b6
          21431 => x"80", -- $053b7
          21432 => x"80", -- $053b8
          21433 => x"80", -- $053b9
          21434 => x"80", -- $053ba
          21435 => x"80", -- $053bb
          21436 => x"80", -- $053bc
          21437 => x"80", -- $053bd
          21438 => x"80", -- $053be
          21439 => x"80", -- $053bf
          21440 => x"80", -- $053c0
          21441 => x"80", -- $053c1
          21442 => x"80", -- $053c2
          21443 => x"80", -- $053c3
          21444 => x"80", -- $053c4
          21445 => x"80", -- $053c5
          21446 => x"80", -- $053c6
          21447 => x"80", -- $053c7
          21448 => x"80", -- $053c8
          21449 => x"80", -- $053c9
          21450 => x"80", -- $053ca
          21451 => x"80", -- $053cb
          21452 => x"80", -- $053cc
          21453 => x"80", -- $053cd
          21454 => x"80", -- $053ce
          21455 => x"80", -- $053cf
          21456 => x"80", -- $053d0
          21457 => x"80", -- $053d1
          21458 => x"80", -- $053d2
          21459 => x"80", -- $053d3
          21460 => x"80", -- $053d4
          21461 => x"80", -- $053d5
          21462 => x"80", -- $053d6
          21463 => x"80", -- $053d7
          21464 => x"80", -- $053d8
          21465 => x"80", -- $053d9
          21466 => x"80", -- $053da
          21467 => x"80", -- $053db
          21468 => x"80", -- $053dc
          21469 => x"80", -- $053dd
          21470 => x"80", -- $053de
          21471 => x"80", -- $053df
          21472 => x"80", -- $053e0
          21473 => x"81", -- $053e1
          21474 => x"81", -- $053e2
          21475 => x"81", -- $053e3
          21476 => x"81", -- $053e4
          21477 => x"81", -- $053e5
          21478 => x"81", -- $053e6
          21479 => x"81", -- $053e7
          21480 => x"81", -- $053e8
          21481 => x"82", -- $053e9
          21482 => x"82", -- $053ea
          21483 => x"82", -- $053eb
          21484 => x"82", -- $053ec
          21485 => x"82", -- $053ed
          21486 => x"82", -- $053ee
          21487 => x"82", -- $053ef
          21488 => x"82", -- $053f0
          21489 => x"82", -- $053f1
          21490 => x"81", -- $053f2
          21491 => x"81", -- $053f3
          21492 => x"81", -- $053f4
          21493 => x"81", -- $053f5
          21494 => x"81", -- $053f6
          21495 => x"81", -- $053f7
          21496 => x"81", -- $053f8
          21497 => x"81", -- $053f9
          21498 => x"81", -- $053fa
          21499 => x"81", -- $053fb
          21500 => x"81", -- $053fc
          21501 => x"81", -- $053fd
          21502 => x"81", -- $053fe
          21503 => x"81", -- $053ff
          21504 => x"81", -- $05400
          21505 => x"81", -- $05401
          21506 => x"81", -- $05402
          21507 => x"80", -- $05403
          21508 => x"80", -- $05404
          21509 => x"80", -- $05405
          21510 => x"80", -- $05406
          21511 => x"81", -- $05407
          21512 => x"81", -- $05408
          21513 => x"81", -- $05409
          21514 => x"81", -- $0540a
          21515 => x"81", -- $0540b
          21516 => x"81", -- $0540c
          21517 => x"81", -- $0540d
          21518 => x"81", -- $0540e
          21519 => x"81", -- $0540f
          21520 => x"81", -- $05410
          21521 => x"81", -- $05411
          21522 => x"81", -- $05412
          21523 => x"81", -- $05413
          21524 => x"81", -- $05414
          21525 => x"81", -- $05415
          21526 => x"81", -- $05416
          21527 => x"81", -- $05417
          21528 => x"80", -- $05418
          21529 => x"80", -- $05419
          21530 => x"81", -- $0541a
          21531 => x"80", -- $0541b
          21532 => x"80", -- $0541c
          21533 => x"81", -- $0541d
          21534 => x"81", -- $0541e
          21535 => x"81", -- $0541f
          21536 => x"81", -- $05420
          21537 => x"81", -- $05421
          21538 => x"81", -- $05422
          21539 => x"81", -- $05423
          21540 => x"81", -- $05424
          21541 => x"81", -- $05425
          21542 => x"82", -- $05426
          21543 => x"81", -- $05427
          21544 => x"81", -- $05428
          21545 => x"81", -- $05429
          21546 => x"82", -- $0542a
          21547 => x"81", -- $0542b
          21548 => x"82", -- $0542c
          21549 => x"82", -- $0542d
          21550 => x"82", -- $0542e
          21551 => x"82", -- $0542f
          21552 => x"82", -- $05430
          21553 => x"82", -- $05431
          21554 => x"82", -- $05432
          21555 => x"82", -- $05433
          21556 => x"82", -- $05434
          21557 => x"82", -- $05435
          21558 => x"82", -- $05436
          21559 => x"82", -- $05437
          21560 => x"82", -- $05438
          21561 => x"82", -- $05439
          21562 => x"81", -- $0543a
          21563 => x"81", -- $0543b
          21564 => x"81", -- $0543c
          21565 => x"81", -- $0543d
          21566 => x"81", -- $0543e
          21567 => x"81", -- $0543f
          21568 => x"81", -- $05440
          21569 => x"81", -- $05441
          21570 => x"81", -- $05442
          21571 => x"80", -- $05443
          21572 => x"80", -- $05444
          21573 => x"80", -- $05445
          21574 => x"80", -- $05446
          21575 => x"80", -- $05447
          21576 => x"80", -- $05448
          21577 => x"80", -- $05449
          21578 => x"80", -- $0544a
          21579 => x"80", -- $0544b
          21580 => x"80", -- $0544c
          21581 => x"80", -- $0544d
          21582 => x"80", -- $0544e
          21583 => x"81", -- $0544f
          21584 => x"81", -- $05450
          21585 => x"81", -- $05451
          21586 => x"81", -- $05452
          21587 => x"81", -- $05453
          21588 => x"81", -- $05454
          21589 => x"81", -- $05455
          21590 => x"81", -- $05456
          21591 => x"82", -- $05457
          21592 => x"82", -- $05458
          21593 => x"82", -- $05459
          21594 => x"82", -- $0545a
          21595 => x"82", -- $0545b
          21596 => x"82", -- $0545c
          21597 => x"82", -- $0545d
          21598 => x"82", -- $0545e
          21599 => x"82", -- $0545f
          21600 => x"82", -- $05460
          21601 => x"82", -- $05461
          21602 => x"82", -- $05462
          21603 => x"82", -- $05463
          21604 => x"82", -- $05464
          21605 => x"82", -- $05465
          21606 => x"82", -- $05466
          21607 => x"82", -- $05467
          21608 => x"82", -- $05468
          21609 => x"82", -- $05469
          21610 => x"82", -- $0546a
          21611 => x"82", -- $0546b
          21612 => x"81", -- $0546c
          21613 => x"81", -- $0546d
          21614 => x"82", -- $0546e
          21615 => x"82", -- $0546f
          21616 => x"82", -- $05470
          21617 => x"82", -- $05471
          21618 => x"82", -- $05472
          21619 => x"82", -- $05473
          21620 => x"82", -- $05474
          21621 => x"82", -- $05475
          21622 => x"82", -- $05476
          21623 => x"82", -- $05477
          21624 => x"82", -- $05478
          21625 => x"82", -- $05479
          21626 => x"82", -- $0547a
          21627 => x"81", -- $0547b
          21628 => x"81", -- $0547c
          21629 => x"81", -- $0547d
          21630 => x"81", -- $0547e
          21631 => x"81", -- $0547f
          21632 => x"81", -- $05480
          21633 => x"81", -- $05481
          21634 => x"81", -- $05482
          21635 => x"81", -- $05483
          21636 => x"81", -- $05484
          21637 => x"81", -- $05485
          21638 => x"81", -- $05486
          21639 => x"81", -- $05487
          21640 => x"81", -- $05488
          21641 => x"81", -- $05489
          21642 => x"80", -- $0548a
          21643 => x"81", -- $0548b
          21644 => x"81", -- $0548c
          21645 => x"81", -- $0548d
          21646 => x"81", -- $0548e
          21647 => x"81", -- $0548f
          21648 => x"80", -- $05490
          21649 => x"80", -- $05491
          21650 => x"80", -- $05492
          21651 => x"80", -- $05493
          21652 => x"80", -- $05494
          21653 => x"80", -- $05495
          21654 => x"81", -- $05496
          21655 => x"81", -- $05497
          21656 => x"81", -- $05498
          21657 => x"81", -- $05499
          21658 => x"81", -- $0549a
          21659 => x"81", -- $0549b
          21660 => x"81", -- $0549c
          21661 => x"81", -- $0549d
          21662 => x"81", -- $0549e
          21663 => x"81", -- $0549f
          21664 => x"82", -- $054a0
          21665 => x"82", -- $054a1
          21666 => x"82", -- $054a2
          21667 => x"82", -- $054a3
          21668 => x"82", -- $054a4
          21669 => x"82", -- $054a5
          21670 => x"82", -- $054a6
          21671 => x"82", -- $054a7
          21672 => x"82", -- $054a8
          21673 => x"81", -- $054a9
          21674 => x"81", -- $054aa
          21675 => x"81", -- $054ab
          21676 => x"81", -- $054ac
          21677 => x"81", -- $054ad
          21678 => x"81", -- $054ae
          21679 => x"81", -- $054af
          21680 => x"81", -- $054b0
          21681 => x"81", -- $054b1
          21682 => x"81", -- $054b2
          21683 => x"81", -- $054b3
          21684 => x"81", -- $054b4
          21685 => x"81", -- $054b5
          21686 => x"81", -- $054b6
          21687 => x"81", -- $054b7
          21688 => x"81", -- $054b8
          21689 => x"81", -- $054b9
          21690 => x"81", -- $054ba
          21691 => x"81", -- $054bb
          21692 => x"81", -- $054bc
          21693 => x"81", -- $054bd
          21694 => x"81", -- $054be
          21695 => x"81", -- $054bf
          21696 => x"81", -- $054c0
          21697 => x"81", -- $054c1
          21698 => x"80", -- $054c2
          21699 => x"80", -- $054c3
          21700 => x"80", -- $054c4
          21701 => x"81", -- $054c5
          21702 => x"81", -- $054c6
          21703 => x"81", -- $054c7
          21704 => x"81", -- $054c8
          21705 => x"81", -- $054c9
          21706 => x"81", -- $054ca
          21707 => x"81", -- $054cb
          21708 => x"81", -- $054cc
          21709 => x"81", -- $054cd
          21710 => x"81", -- $054ce
          21711 => x"81", -- $054cf
          21712 => x"81", -- $054d0
          21713 => x"81", -- $054d1
          21714 => x"81", -- $054d2
          21715 => x"81", -- $054d3
          21716 => x"81", -- $054d4
          21717 => x"81", -- $054d5
          21718 => x"81", -- $054d6
          21719 => x"81", -- $054d7
          21720 => x"81", -- $054d8
          21721 => x"81", -- $054d9
          21722 => x"81", -- $054da
          21723 => x"81", -- $054db
          21724 => x"81", -- $054dc
          21725 => x"81", -- $054dd
          21726 => x"81", -- $054de
          21727 => x"81", -- $054df
          21728 => x"81", -- $054e0
          21729 => x"80", -- $054e1
          21730 => x"80", -- $054e2
          21731 => x"80", -- $054e3
          21732 => x"80", -- $054e4
          21733 => x"80", -- $054e5
          21734 => x"80", -- $054e6
          21735 => x"81", -- $054e7
          21736 => x"81", -- $054e8
          21737 => x"80", -- $054e9
          21738 => x"80", -- $054ea
          21739 => x"80", -- $054eb
          21740 => x"80", -- $054ec
          21741 => x"80", -- $054ed
          21742 => x"80", -- $054ee
          21743 => x"80", -- $054ef
          21744 => x"80", -- $054f0
          21745 => x"80", -- $054f1
          21746 => x"81", -- $054f2
          21747 => x"81", -- $054f3
          21748 => x"81", -- $054f4
          21749 => x"81", -- $054f5
          21750 => x"81", -- $054f6
          21751 => x"81", -- $054f7
          21752 => x"81", -- $054f8
          21753 => x"81", -- $054f9
          21754 => x"81", -- $054fa
          21755 => x"80", -- $054fb
          21756 => x"80", -- $054fc
          21757 => x"80", -- $054fd
          21758 => x"80", -- $054fe
          21759 => x"80", -- $054ff
          21760 => x"80", -- $05500
          21761 => x"80", -- $05501
          21762 => x"80", -- $05502
          21763 => x"80", -- $05503
          21764 => x"80", -- $05504
          21765 => x"80", -- $05505
          21766 => x"80", -- $05506
          21767 => x"80", -- $05507
          21768 => x"80", -- $05508
          21769 => x"80", -- $05509
          21770 => x"80", -- $0550a
          21771 => x"80", -- $0550b
          21772 => x"80", -- $0550c
          21773 => x"80", -- $0550d
          21774 => x"80", -- $0550e
          21775 => x"80", -- $0550f
          21776 => x"80", -- $05510
          21777 => x"80", -- $05511
          21778 => x"80", -- $05512
          21779 => x"80", -- $05513
          21780 => x"80", -- $05514
          21781 => x"80", -- $05515
          21782 => x"80", -- $05516
          21783 => x"80", -- $05517
          21784 => x"80", -- $05518
          21785 => x"80", -- $05519
          21786 => x"80", -- $0551a
          21787 => x"81", -- $0551b
          21788 => x"81", -- $0551c
          21789 => x"81", -- $0551d
          21790 => x"81", -- $0551e
          21791 => x"81", -- $0551f
          21792 => x"81", -- $05520
          21793 => x"81", -- $05521
          21794 => x"81", -- $05522
          21795 => x"81", -- $05523
          21796 => x"80", -- $05524
          21797 => x"80", -- $05525
          21798 => x"80", -- $05526
          21799 => x"80", -- $05527
          21800 => x"80", -- $05528
          21801 => x"80", -- $05529
          21802 => x"80", -- $0552a
          21803 => x"80", -- $0552b
          21804 => x"80", -- $0552c
          21805 => x"80", -- $0552d
          21806 => x"80", -- $0552e
          21807 => x"80", -- $0552f
          21808 => x"80", -- $05530
          21809 => x"80", -- $05531
          21810 => x"80", -- $05532
          21811 => x"80", -- $05533
          21812 => x"80", -- $05534
          21813 => x"80", -- $05535
          21814 => x"80", -- $05536
          21815 => x"80", -- $05537
          21816 => x"80", -- $05538
          21817 => x"80", -- $05539
          21818 => x"80", -- $0553a
          21819 => x"80", -- $0553b
          21820 => x"80", -- $0553c
          21821 => x"80", -- $0553d
          21822 => x"80", -- $0553e
          21823 => x"80", -- $0553f
          21824 => x"80", -- $05540
          21825 => x"80", -- $05541
          21826 => x"80", -- $05542
          21827 => x"80", -- $05543
          21828 => x"80", -- $05544
          21829 => x"80", -- $05545
          21830 => x"80", -- $05546
          21831 => x"80", -- $05547
          21832 => x"80", -- $05548
          21833 => x"80", -- $05549
          21834 => x"80", -- $0554a
          21835 => x"7f", -- $0554b
          21836 => x"80", -- $0554c
          21837 => x"80", -- $0554d
          21838 => x"80", -- $0554e
          21839 => x"80", -- $0554f
          21840 => x"80", -- $05550
          21841 => x"80", -- $05551
          21842 => x"80", -- $05552
          21843 => x"80", -- $05553
          21844 => x"80", -- $05554
          21845 => x"80", -- $05555
          21846 => x"80", -- $05556
          21847 => x"80", -- $05557
          21848 => x"80", -- $05558
          21849 => x"80", -- $05559
          21850 => x"80", -- $0555a
          21851 => x"80", -- $0555b
          21852 => x"80", -- $0555c
          21853 => x"80", -- $0555d
          21854 => x"80", -- $0555e
          21855 => x"80", -- $0555f
          21856 => x"80", -- $05560
          21857 => x"7f", -- $05561
          21858 => x"7f", -- $05562
          21859 => x"7f", -- $05563
          21860 => x"7f", -- $05564
          21861 => x"7f", -- $05565
          21862 => x"7f", -- $05566
          21863 => x"7f", -- $05567
          21864 => x"7f", -- $05568
          21865 => x"7f", -- $05569
          21866 => x"7f", -- $0556a
          21867 => x"7f", -- $0556b
          21868 => x"7f", -- $0556c
          21869 => x"7f", -- $0556d
          21870 => x"7f", -- $0556e
          21871 => x"7f", -- $0556f
          21872 => x"7f", -- $05570
          21873 => x"7f", -- $05571
          21874 => x"7f", -- $05572
          21875 => x"7f", -- $05573
          21876 => x"7f", -- $05574
          21877 => x"7f", -- $05575
          21878 => x"7f", -- $05576
          21879 => x"7f", -- $05577
          21880 => x"7f", -- $05578
          21881 => x"7f", -- $05579
          21882 => x"7f", -- $0557a
          21883 => x"7f", -- $0557b
          21884 => x"7f", -- $0557c
          21885 => x"7f", -- $0557d
          21886 => x"7e", -- $0557e
          21887 => x"7e", -- $0557f
          21888 => x"7e", -- $05580
          21889 => x"7e", -- $05581
          21890 => x"7e", -- $05582
          21891 => x"7e", -- $05583
          21892 => x"7e", -- $05584
          21893 => x"7e", -- $05585
          21894 => x"7e", -- $05586
          21895 => x"7e", -- $05587
          21896 => x"7f", -- $05588
          21897 => x"7f", -- $05589
          21898 => x"7e", -- $0558a
          21899 => x"7f", -- $0558b
          21900 => x"7f", -- $0558c
          21901 => x"7f", -- $0558d
          21902 => x"7f", -- $0558e
          21903 => x"7f", -- $0558f
          21904 => x"7f", -- $05590
          21905 => x"7f", -- $05591
          21906 => x"7f", -- $05592
          21907 => x"7f", -- $05593
          21908 => x"7f", -- $05594
          21909 => x"7f", -- $05595
          21910 => x"7f", -- $05596
          21911 => x"7f", -- $05597
          21912 => x"7f", -- $05598
          21913 => x"7f", -- $05599
          21914 => x"7f", -- $0559a
          21915 => x"7f", -- $0559b
          21916 => x"7f", -- $0559c
          21917 => x"7f", -- $0559d
          21918 => x"7f", -- $0559e
          21919 => x"7f", -- $0559f
          21920 => x"7f", -- $055a0
          21921 => x"7f", -- $055a1
          21922 => x"7f", -- $055a2
          21923 => x"7e", -- $055a3
          21924 => x"7e", -- $055a4
          21925 => x"7e", -- $055a5
          21926 => x"7e", -- $055a6
          21927 => x"7e", -- $055a7
          21928 => x"7f", -- $055a8
          21929 => x"7f", -- $055a9
          21930 => x"7f", -- $055aa
          21931 => x"7f", -- $055ab
          21932 => x"7f", -- $055ac
          21933 => x"7f", -- $055ad
          21934 => x"7f", -- $055ae
          21935 => x"7f", -- $055af
          21936 => x"7f", -- $055b0
          21937 => x"7f", -- $055b1
          21938 => x"7f", -- $055b2
          21939 => x"7f", -- $055b3
          21940 => x"7f", -- $055b4
          21941 => x"7f", -- $055b5
          21942 => x"7f", -- $055b6
          21943 => x"7f", -- $055b7
          21944 => x"7f", -- $055b8
          21945 => x"7f", -- $055b9
          21946 => x"7f", -- $055ba
          21947 => x"7f", -- $055bb
          21948 => x"7f", -- $055bc
          21949 => x"7f", -- $055bd
          21950 => x"7f", -- $055be
          21951 => x"7f", -- $055bf
          21952 => x"7f", -- $055c0
          21953 => x"7f", -- $055c1
          21954 => x"7f", -- $055c2
          21955 => x"7f", -- $055c3
          21956 => x"7f", -- $055c4
          21957 => x"7f", -- $055c5
          21958 => x"7f", -- $055c6
          21959 => x"7f", -- $055c7
          21960 => x"7f", -- $055c8
          21961 => x"7f", -- $055c9
          21962 => x"7f", -- $055ca
          21963 => x"7f", -- $055cb
          21964 => x"7f", -- $055cc
          21965 => x"7f", -- $055cd
          21966 => x"7f", -- $055ce
          21967 => x"7f", -- $055cf
          21968 => x"7f", -- $055d0
          21969 => x"7f", -- $055d1
          21970 => x"80", -- $055d2
          21971 => x"80", -- $055d3
          21972 => x"80", -- $055d4
          21973 => x"80", -- $055d5
          21974 => x"80", -- $055d6
          21975 => x"7f", -- $055d7
          21976 => x"7f", -- $055d8
          21977 => x"7f", -- $055d9
          21978 => x"7f", -- $055da
          21979 => x"7f", -- $055db
          21980 => x"7f", -- $055dc
          21981 => x"7f", -- $055dd
          21982 => x"7f", -- $055de
          21983 => x"7f", -- $055df
          21984 => x"7f", -- $055e0
          21985 => x"7f", -- $055e1
          21986 => x"7f", -- $055e2
          21987 => x"7f", -- $055e3
          21988 => x"7f", -- $055e4
          21989 => x"7f", -- $055e5
          21990 => x"7f", -- $055e6
          21991 => x"7f", -- $055e7
          21992 => x"7f", -- $055e8
          21993 => x"7f", -- $055e9
          21994 => x"7f", -- $055ea
          21995 => x"7f", -- $055eb
          21996 => x"7f", -- $055ec
          21997 => x"7f", -- $055ed
          21998 => x"7f", -- $055ee
          21999 => x"7f", -- $055ef
          22000 => x"7f", -- $055f0
          22001 => x"7f", -- $055f1
          22002 => x"7f", -- $055f2
          22003 => x"7f", -- $055f3
          22004 => x"7f", -- $055f4
          22005 => x"7f", -- $055f5
          22006 => x"7f", -- $055f6
          22007 => x"7f", -- $055f7
          22008 => x"7f", -- $055f8
          22009 => x"7f", -- $055f9
          22010 => x"7f", -- $055fa
          22011 => x"7f", -- $055fb
          22012 => x"7f", -- $055fc
          22013 => x"7f", -- $055fd
          22014 => x"7f", -- $055fe
          22015 => x"7f", -- $055ff
          22016 => x"7f", -- $05600
          22017 => x"7f", -- $05601
          22018 => x"7f", -- $05602
          22019 => x"7f", -- $05603
          22020 => x"7f", -- $05604
          22021 => x"7f", -- $05605
          22022 => x"7f", -- $05606
          22023 => x"7f", -- $05607
          22024 => x"7f", -- $05608
          22025 => x"7f", -- $05609
          22026 => x"7f", -- $0560a
          22027 => x"7f", -- $0560b
          22028 => x"7f", -- $0560c
          22029 => x"7f", -- $0560d
          22030 => x"7f", -- $0560e
          22031 => x"7f", -- $0560f
          22032 => x"7f", -- $05610
          22033 => x"7f", -- $05611
          22034 => x"7f", -- $05612
          22035 => x"7f", -- $05613
          22036 => x"7f", -- $05614
          22037 => x"7f", -- $05615
          22038 => x"7f", -- $05616
          22039 => x"7f", -- $05617
          22040 => x"7f", -- $05618
          22041 => x"7f", -- $05619
          22042 => x"7f", -- $0561a
          22043 => x"7f", -- $0561b
          22044 => x"7f", -- $0561c
          22045 => x"7f", -- $0561d
          22046 => x"7f", -- $0561e
          22047 => x"7e", -- $0561f
          22048 => x"7e", -- $05620
          22049 => x"7e", -- $05621
          22050 => x"7e", -- $05622
          22051 => x"7f", -- $05623
          22052 => x"7f", -- $05624
          22053 => x"7e", -- $05625
          22054 => x"7e", -- $05626
          22055 => x"7e", -- $05627
          22056 => x"7e", -- $05628
          22057 => x"7f", -- $05629
          22058 => x"7f", -- $0562a
          22059 => x"7f", -- $0562b
          22060 => x"7f", -- $0562c
          22061 => x"7f", -- $0562d
          22062 => x"7f", -- $0562e
          22063 => x"7f", -- $0562f
          22064 => x"7f", -- $05630
          22065 => x"7f", -- $05631
          22066 => x"7f", -- $05632
          22067 => x"7f", -- $05633
          22068 => x"7f", -- $05634
          22069 => x"7e", -- $05635
          22070 => x"7e", -- $05636
          22071 => x"7e", -- $05637
          22072 => x"7e", -- $05638
          22073 => x"7f", -- $05639
          22074 => x"7f", -- $0563a
          22075 => x"7f", -- $0563b
          22076 => x"7f", -- $0563c
          22077 => x"7f", -- $0563d
          22078 => x"7f", -- $0563e
          22079 => x"7f", -- $0563f
          22080 => x"7e", -- $05640
          22081 => x"7f", -- $05641
          22082 => x"7e", -- $05642
          22083 => x"7f", -- $05643
          22084 => x"7f", -- $05644
          22085 => x"7f", -- $05645
          22086 => x"7f", -- $05646
          22087 => x"7f", -- $05647
          22088 => x"7f", -- $05648
          22089 => x"7f", -- $05649
          22090 => x"7f", -- $0564a
          22091 => x"7f", -- $0564b
          22092 => x"7f", -- $0564c
          22093 => x"7f", -- $0564d
          22094 => x"7f", -- $0564e
          22095 => x"7f", -- $0564f
          22096 => x"7f", -- $05650
          22097 => x"7f", -- $05651
          22098 => x"7f", -- $05652
          22099 => x"7f", -- $05653
          22100 => x"7f", -- $05654
          22101 => x"7f", -- $05655
          22102 => x"7f", -- $05656
          22103 => x"7f", -- $05657
          22104 => x"7f", -- $05658
          22105 => x"7f", -- $05659
          22106 => x"7f", -- $0565a
          22107 => x"7f", -- $0565b
          22108 => x"7f", -- $0565c
          22109 => x"7f", -- $0565d
          22110 => x"7f", -- $0565e
          22111 => x"7f", -- $0565f
          22112 => x"7f", -- $05660
          22113 => x"7f", -- $05661
          22114 => x"80", -- $05662
          22115 => x"80", -- $05663
          22116 => x"80", -- $05664
          22117 => x"7f", -- $05665
          22118 => x"7f", -- $05666
          22119 => x"7f", -- $05667
          22120 => x"80", -- $05668
          22121 => x"80", -- $05669
          22122 => x"80", -- $0566a
          22123 => x"80", -- $0566b
          22124 => x"80", -- $0566c
          22125 => x"80", -- $0566d
          22126 => x"80", -- $0566e
          22127 => x"80", -- $0566f
          22128 => x"80", -- $05670
          22129 => x"80", -- $05671
          22130 => x"80", -- $05672
          22131 => x"80", -- $05673
          22132 => x"80", -- $05674
          22133 => x"80", -- $05675
          22134 => x"80", -- $05676
          22135 => x"80", -- $05677
          22136 => x"80", -- $05678
          22137 => x"80", -- $05679
          22138 => x"80", -- $0567a
          22139 => x"80", -- $0567b
          22140 => x"80", -- $0567c
          22141 => x"80", -- $0567d
          22142 => x"80", -- $0567e
          22143 => x"80", -- $0567f
          22144 => x"80", -- $05680
          22145 => x"80", -- $05681
          22146 => x"80", -- $05682
          22147 => x"80", -- $05683
          22148 => x"80", -- $05684
          22149 => x"80", -- $05685
          22150 => x"80", -- $05686
          22151 => x"80", -- $05687
          22152 => x"80", -- $05688
          22153 => x"80", -- $05689
          22154 => x"80", -- $0568a
          22155 => x"80", -- $0568b
          22156 => x"80", -- $0568c
          22157 => x"80", -- $0568d
          22158 => x"80", -- $0568e
          22159 => x"80", -- $0568f
          22160 => x"80", -- $05690
          22161 => x"80", -- $05691
          22162 => x"80", -- $05692
          22163 => x"80", -- $05693
          22164 => x"80", -- $05694
          22165 => x"80", -- $05695
          22166 => x"80", -- $05696
          22167 => x"80", -- $05697
          22168 => x"80", -- $05698
          22169 => x"80", -- $05699
          22170 => x"80", -- $0569a
          22171 => x"80", -- $0569b
          22172 => x"80", -- $0569c
          22173 => x"80", -- $0569d
          22174 => x"80", -- $0569e
          22175 => x"80", -- $0569f
          22176 => x"80", -- $056a0
          22177 => x"80", -- $056a1
          22178 => x"80", -- $056a2
          22179 => x"80", -- $056a3
          22180 => x"80", -- $056a4
          22181 => x"80", -- $056a5
          22182 => x"80", -- $056a6
          22183 => x"80", -- $056a7
          22184 => x"80", -- $056a8
          22185 => x"80", -- $056a9
          22186 => x"80", -- $056aa
          22187 => x"80", -- $056ab
          22188 => x"80", -- $056ac
          22189 => x"80", -- $056ad
          22190 => x"80", -- $056ae
          22191 => x"80", -- $056af
          22192 => x"80", -- $056b0
          22193 => x"80", -- $056b1
          22194 => x"80", -- $056b2
          22195 => x"80", -- $056b3
          22196 => x"80", -- $056b4
          22197 => x"80", -- $056b5
          22198 => x"80", -- $056b6
          22199 => x"81", -- $056b7
          22200 => x"81", -- $056b8
          22201 => x"81", -- $056b9
          22202 => x"81", -- $056ba
          22203 => x"81", -- $056bb
          22204 => x"81", -- $056bc
          22205 => x"81", -- $056bd
          22206 => x"81", -- $056be
          22207 => x"81", -- $056bf
          22208 => x"81", -- $056c0
          22209 => x"81", -- $056c1
          22210 => x"81", -- $056c2
          22211 => x"81", -- $056c3
          22212 => x"81", -- $056c4
          22213 => x"81", -- $056c5
          22214 => x"81", -- $056c6
          22215 => x"81", -- $056c7
          22216 => x"81", -- $056c8
          22217 => x"81", -- $056c9
          22218 => x"81", -- $056ca
          22219 => x"81", -- $056cb
          22220 => x"81", -- $056cc
          22221 => x"81", -- $056cd
          22222 => x"81", -- $056ce
          22223 => x"81", -- $056cf
          22224 => x"81", -- $056d0
          22225 => x"81", -- $056d1
          22226 => x"81", -- $056d2
          22227 => x"81", -- $056d3
          22228 => x"81", -- $056d4
          22229 => x"81", -- $056d5
          22230 => x"81", -- $056d6
          22231 => x"81", -- $056d7
          22232 => x"81", -- $056d8
          22233 => x"81", -- $056d9
          22234 => x"81", -- $056da
          22235 => x"81", -- $056db
          22236 => x"81", -- $056dc
          22237 => x"81", -- $056dd
          22238 => x"81", -- $056de
          22239 => x"81", -- $056df
          22240 => x"81", -- $056e0
          22241 => x"81", -- $056e1
          22242 => x"81", -- $056e2
          22243 => x"81", -- $056e3
          22244 => x"81", -- $056e4
          22245 => x"81", -- $056e5
          22246 => x"81", -- $056e6
          22247 => x"81", -- $056e7
          22248 => x"81", -- $056e8
          22249 => x"81", -- $056e9
          22250 => x"81", -- $056ea
          22251 => x"81", -- $056eb
          22252 => x"81", -- $056ec
          22253 => x"81", -- $056ed
          22254 => x"81", -- $056ee
          22255 => x"81", -- $056ef
          22256 => x"81", -- $056f0
          22257 => x"81", -- $056f1
          22258 => x"81", -- $056f2
          22259 => x"81", -- $056f3
          22260 => x"81", -- $056f4
          22261 => x"81", -- $056f5
          22262 => x"81", -- $056f6
          22263 => x"81", -- $056f7
          22264 => x"81", -- $056f8
          22265 => x"81", -- $056f9
          22266 => x"81", -- $056fa
          22267 => x"81", -- $056fb
          22268 => x"81", -- $056fc
          22269 => x"81", -- $056fd
          22270 => x"81", -- $056fe
          22271 => x"81", -- $056ff
          22272 => x"81", -- $05700
          22273 => x"81", -- $05701
          22274 => x"81", -- $05702
          22275 => x"81", -- $05703
          22276 => x"81", -- $05704
          22277 => x"81", -- $05705
          22278 => x"81", -- $05706
          22279 => x"81", -- $05707
          22280 => x"81", -- $05708
          22281 => x"81", -- $05709
          22282 => x"81", -- $0570a
          22283 => x"81", -- $0570b
          22284 => x"81", -- $0570c
          22285 => x"81", -- $0570d
          22286 => x"81", -- $0570e
          22287 => x"81", -- $0570f
          22288 => x"82", -- $05710
          22289 => x"82", -- $05711
          22290 => x"81", -- $05712
          22291 => x"81", -- $05713
          22292 => x"81", -- $05714
          22293 => x"81", -- $05715
          22294 => x"81", -- $05716
          22295 => x"81", -- $05717
          22296 => x"81", -- $05718
          22297 => x"81", -- $05719
          22298 => x"81", -- $0571a
          22299 => x"81", -- $0571b
          22300 => x"81", -- $0571c
          22301 => x"81", -- $0571d
          22302 => x"81", -- $0571e
          22303 => x"81", -- $0571f
          22304 => x"81", -- $05720
          22305 => x"81", -- $05721
          22306 => x"81", -- $05722
          22307 => x"81", -- $05723
          22308 => x"81", -- $05724
          22309 => x"81", -- $05725
          22310 => x"81", -- $05726
          22311 => x"81", -- $05727
          22312 => x"81", -- $05728
          22313 => x"81", -- $05729
          22314 => x"81", -- $0572a
          22315 => x"81", -- $0572b
          22316 => x"81", -- $0572c
          22317 => x"81", -- $0572d
          22318 => x"81", -- $0572e
          22319 => x"81", -- $0572f
          22320 => x"81", -- $05730
          22321 => x"81", -- $05731
          22322 => x"81", -- $05732
          22323 => x"81", -- $05733
          22324 => x"81", -- $05734
          22325 => x"81", -- $05735
          22326 => x"81", -- $05736
          22327 => x"81", -- $05737
          22328 => x"81", -- $05738
          22329 => x"81", -- $05739
          22330 => x"81", -- $0573a
          22331 => x"81", -- $0573b
          22332 => x"81", -- $0573c
          22333 => x"81", -- $0573d
          22334 => x"81", -- $0573e
          22335 => x"81", -- $0573f
          22336 => x"81", -- $05740
          22337 => x"81", -- $05741
          22338 => x"80", -- $05742
          22339 => x"80", -- $05743
          22340 => x"80", -- $05744
          22341 => x"80", -- $05745
          22342 => x"80", -- $05746
          22343 => x"80", -- $05747
          22344 => x"80", -- $05748
          22345 => x"80", -- $05749
          22346 => x"80", -- $0574a
          22347 => x"80", -- $0574b
          22348 => x"80", -- $0574c
          22349 => x"81", -- $0574d
          22350 => x"81", -- $0574e
          22351 => x"81", -- $0574f
          22352 => x"81", -- $05750
          22353 => x"81", -- $05751
          22354 => x"81", -- $05752
          22355 => x"81", -- $05753
          22356 => x"81", -- $05754
          22357 => x"81", -- $05755
          22358 => x"81", -- $05756
          22359 => x"81", -- $05757
          22360 => x"81", -- $05758
          22361 => x"81", -- $05759
          22362 => x"81", -- $0575a
          22363 => x"80", -- $0575b
          22364 => x"81", -- $0575c
          22365 => x"81", -- $0575d
          22366 => x"81", -- $0575e
          22367 => x"81", -- $0575f
          22368 => x"81", -- $05760
          22369 => x"81", -- $05761
          22370 => x"81", -- $05762
          22371 => x"81", -- $05763
          22372 => x"81", -- $05764
          22373 => x"81", -- $05765
          22374 => x"81", -- $05766
          22375 => x"81", -- $05767
          22376 => x"81", -- $05768
          22377 => x"81", -- $05769
          22378 => x"81", -- $0576a
          22379 => x"81", -- $0576b
          22380 => x"81", -- $0576c
          22381 => x"81", -- $0576d
          22382 => x"81", -- $0576e
          22383 => x"81", -- $0576f
          22384 => x"81", -- $05770
          22385 => x"81", -- $05771
          22386 => x"82", -- $05772
          22387 => x"82", -- $05773
          22388 => x"82", -- $05774
          22389 => x"82", -- $05775
          22390 => x"82", -- $05776
          22391 => x"82", -- $05777
          22392 => x"82", -- $05778
          22393 => x"82", -- $05779
          22394 => x"82", -- $0577a
          22395 => x"82", -- $0577b
          22396 => x"82", -- $0577c
          22397 => x"82", -- $0577d
          22398 => x"82", -- $0577e
          22399 => x"82", -- $0577f
          22400 => x"82", -- $05780
          22401 => x"82", -- $05781
          22402 => x"82", -- $05782
          22403 => x"82", -- $05783
          22404 => x"82", -- $05784
          22405 => x"82", -- $05785
          22406 => x"82", -- $05786
          22407 => x"82", -- $05787
          22408 => x"82", -- $05788
          22409 => x"82", -- $05789
          22410 => x"82", -- $0578a
          22411 => x"82", -- $0578b
          22412 => x"82", -- $0578c
          22413 => x"82", -- $0578d
          22414 => x"82", -- $0578e
          22415 => x"82", -- $0578f
          22416 => x"82", -- $05790
          22417 => x"82", -- $05791
          22418 => x"82", -- $05792
          22419 => x"82", -- $05793
          22420 => x"82", -- $05794
          22421 => x"82", -- $05795
          22422 => x"82", -- $05796
          22423 => x"82", -- $05797
          22424 => x"82", -- $05798
          22425 => x"82", -- $05799
          22426 => x"82", -- $0579a
          22427 => x"82", -- $0579b
          22428 => x"82", -- $0579c
          22429 => x"82", -- $0579d
          22430 => x"82", -- $0579e
          22431 => x"82", -- $0579f
          22432 => x"82", -- $057a0
          22433 => x"82", -- $057a1
          22434 => x"82", -- $057a2
          22435 => x"82", -- $057a3
          22436 => x"82", -- $057a4
          22437 => x"82", -- $057a5
          22438 => x"82", -- $057a6
          22439 => x"82", -- $057a7
          22440 => x"82", -- $057a8
          22441 => x"82", -- $057a9
          22442 => x"82", -- $057aa
          22443 => x"81", -- $057ab
          22444 => x"81", -- $057ac
          22445 => x"81", -- $057ad
          22446 => x"81", -- $057ae
          22447 => x"81", -- $057af
          22448 => x"81", -- $057b0
          22449 => x"81", -- $057b1
          22450 => x"81", -- $057b2
          22451 => x"81", -- $057b3
          22452 => x"81", -- $057b4
          22453 => x"81", -- $057b5
          22454 => x"81", -- $057b6
          22455 => x"81", -- $057b7
          22456 => x"81", -- $057b8
          22457 => x"81", -- $057b9
          22458 => x"81", -- $057ba
          22459 => x"81", -- $057bb
          22460 => x"81", -- $057bc
          22461 => x"81", -- $057bd
          22462 => x"81", -- $057be
          22463 => x"80", -- $057bf
          22464 => x"80", -- $057c0
          22465 => x"80", -- $057c1
          22466 => x"80", -- $057c2
          22467 => x"80", -- $057c3
          22468 => x"81", -- $057c4
          22469 => x"80", -- $057c5
          22470 => x"80", -- $057c6
          22471 => x"81", -- $057c7
          22472 => x"81", -- $057c8
          22473 => x"80", -- $057c9
          22474 => x"80", -- $057ca
          22475 => x"80", -- $057cb
          22476 => x"80", -- $057cc
          22477 => x"80", -- $057cd
          22478 => x"80", -- $057ce
          22479 => x"80", -- $057cf
          22480 => x"80", -- $057d0
          22481 => x"80", -- $057d1
          22482 => x"80", -- $057d2
          22483 => x"80", -- $057d3
          22484 => x"80", -- $057d4
          22485 => x"80", -- $057d5
          22486 => x"80", -- $057d6
          22487 => x"80", -- $057d7
          22488 => x"80", -- $057d8
          22489 => x"80", -- $057d9
          22490 => x"80", -- $057da
          22491 => x"80", -- $057db
          22492 => x"80", -- $057dc
          22493 => x"80", -- $057dd
          22494 => x"80", -- $057de
          22495 => x"80", -- $057df
          22496 => x"80", -- $057e0
          22497 => x"80", -- $057e1
          22498 => x"80", -- $057e2
          22499 => x"80", -- $057e3
          22500 => x"80", -- $057e4
          22501 => x"80", -- $057e5
          22502 => x"80", -- $057e6
          22503 => x"80", -- $057e7
          22504 => x"80", -- $057e8
          22505 => x"80", -- $057e9
          22506 => x"80", -- $057ea
          22507 => x"80", -- $057eb
          22508 => x"80", -- $057ec
          22509 => x"80", -- $057ed
          22510 => x"80", -- $057ee
          22511 => x"80", -- $057ef
          22512 => x"80", -- $057f0
          22513 => x"80", -- $057f1
          22514 => x"80", -- $057f2
          22515 => x"80", -- $057f3
          22516 => x"80", -- $057f4
          22517 => x"80", -- $057f5
          22518 => x"80", -- $057f6
          22519 => x"80", -- $057f7
          22520 => x"80", -- $057f8
          22521 => x"80", -- $057f9
          22522 => x"80", -- $057fa
          22523 => x"80", -- $057fb
          22524 => x"80", -- $057fc
          22525 => x"80", -- $057fd
          22526 => x"80", -- $057fe
          22527 => x"80", -- $057ff
          22528 => x"7f", -- $05800
          22529 => x"7f", -- $05801
          22530 => x"80", -- $05802
          22531 => x"80", -- $05803
          22532 => x"80", -- $05804
          22533 => x"80", -- $05805
          22534 => x"80", -- $05806
          22535 => x"80", -- $05807
          22536 => x"80", -- $05808
          22537 => x"80", -- $05809
          22538 => x"80", -- $0580a
          22539 => x"80", -- $0580b
          22540 => x"80", -- $0580c
          22541 => x"80", -- $0580d
          22542 => x"80", -- $0580e
          22543 => x"7f", -- $0580f
          22544 => x"7f", -- $05810
          22545 => x"7f", -- $05811
          22546 => x"7f", -- $05812
          22547 => x"7f", -- $05813
          22548 => x"7f", -- $05814
          22549 => x"7f", -- $05815
          22550 => x"7f", -- $05816
          22551 => x"7f", -- $05817
          22552 => x"7f", -- $05818
          22553 => x"7f", -- $05819
          22554 => x"7f", -- $0581a
          22555 => x"7f", -- $0581b
          22556 => x"7f", -- $0581c
          22557 => x"7f", -- $0581d
          22558 => x"7f", -- $0581e
          22559 => x"7f", -- $0581f
          22560 => x"7f", -- $05820
          22561 => x"7f", -- $05821
          22562 => x"7f", -- $05822
          22563 => x"80", -- $05823
          22564 => x"7f", -- $05824
          22565 => x"80", -- $05825
          22566 => x"80", -- $05826
          22567 => x"80", -- $05827
          22568 => x"80", -- $05828
          22569 => x"80", -- $05829
          22570 => x"80", -- $0582a
          22571 => x"80", -- $0582b
          22572 => x"80", -- $0582c
          22573 => x"80", -- $0582d
          22574 => x"80", -- $0582e
          22575 => x"80", -- $0582f
          22576 => x"7f", -- $05830
          22577 => x"7f", -- $05831
          22578 => x"7f", -- $05832
          22579 => x"7f", -- $05833
          22580 => x"7f", -- $05834
          22581 => x"7f", -- $05835
          22582 => x"7f", -- $05836
          22583 => x"7f", -- $05837
          22584 => x"7f", -- $05838
          22585 => x"7f", -- $05839
          22586 => x"7f", -- $0583a
          22587 => x"80", -- $0583b
          22588 => x"80", -- $0583c
          22589 => x"80", -- $0583d
          22590 => x"80", -- $0583e
          22591 => x"80", -- $0583f
          22592 => x"80", -- $05840
          22593 => x"80", -- $05841
          22594 => x"80", -- $05842
          22595 => x"80", -- $05843
          22596 => x"80", -- $05844
          22597 => x"80", -- $05845
          22598 => x"80", -- $05846
          22599 => x"80", -- $05847
          22600 => x"80", -- $05848
          22601 => x"80", -- $05849
          22602 => x"80", -- $0584a
          22603 => x"80", -- $0584b
          22604 => x"80", -- $0584c
          22605 => x"80", -- $0584d
          22606 => x"80", -- $0584e
          22607 => x"80", -- $0584f
          22608 => x"80", -- $05850
          22609 => x"80", -- $05851
          22610 => x"80", -- $05852
          22611 => x"80", -- $05853
          22612 => x"80", -- $05854
          22613 => x"80", -- $05855
          22614 => x"80", -- $05856
          22615 => x"80", -- $05857
          22616 => x"80", -- $05858
          22617 => x"80", -- $05859
          22618 => x"80", -- $0585a
          22619 => x"80", -- $0585b
          22620 => x"80", -- $0585c
          22621 => x"80", -- $0585d
          22622 => x"80", -- $0585e
          22623 => x"80", -- $0585f
          22624 => x"80", -- $05860
          22625 => x"80", -- $05861
          22626 => x"80", -- $05862
          22627 => x"80", -- $05863
          22628 => x"80", -- $05864
          22629 => x"80", -- $05865
          22630 => x"80", -- $05866
          22631 => x"80", -- $05867
          22632 => x"80", -- $05868
          22633 => x"80", -- $05869
          22634 => x"80", -- $0586a
          22635 => x"80", -- $0586b
          22636 => x"80", -- $0586c
          22637 => x"80", -- $0586d
          22638 => x"80", -- $0586e
          22639 => x"80", -- $0586f
          22640 => x"80", -- $05870
          22641 => x"80", -- $05871
          22642 => x"80", -- $05872
          22643 => x"80", -- $05873
          22644 => x"80", -- $05874
          22645 => x"80", -- $05875
          22646 => x"80", -- $05876
          22647 => x"80", -- $05877
          22648 => x"80", -- $05878
          22649 => x"80", -- $05879
          22650 => x"80", -- $0587a
          22651 => x"80", -- $0587b
          22652 => x"80", -- $0587c
          22653 => x"80", -- $0587d
          22654 => x"80", -- $0587e
          22655 => x"80", -- $0587f
          22656 => x"80", -- $05880
          22657 => x"7f", -- $05881
          22658 => x"80", -- $05882
          22659 => x"7f", -- $05883
          22660 => x"7f", -- $05884
          22661 => x"7f", -- $05885
          22662 => x"7f", -- $05886
          22663 => x"7f", -- $05887
          22664 => x"7f", -- $05888
          22665 => x"7f", -- $05889
          22666 => x"7f", -- $0588a
          22667 => x"7f", -- $0588b
          22668 => x"7f", -- $0588c
          22669 => x"7f", -- $0588d
          22670 => x"7f", -- $0588e
          22671 => x"7f", -- $0588f
          22672 => x"7f", -- $05890
          22673 => x"7f", -- $05891
          22674 => x"7f", -- $05892
          22675 => x"80", -- $05893
          22676 => x"80", -- $05894
          22677 => x"80", -- $05895
          22678 => x"80", -- $05896
          22679 => x"7f", -- $05897
          22680 => x"7f", -- $05898
          22681 => x"7f", -- $05899
          22682 => x"7f", -- $0589a
          22683 => x"7f", -- $0589b
          22684 => x"7f", -- $0589c
          22685 => x"7f", -- $0589d
          22686 => x"7f", -- $0589e
          22687 => x"7f", -- $0589f
          22688 => x"7f", -- $058a0
          22689 => x"7f", -- $058a1
          22690 => x"7f", -- $058a2
          22691 => x"7f", -- $058a3
          22692 => x"7f", -- $058a4
          22693 => x"7f", -- $058a5
          22694 => x"7f", -- $058a6
          22695 => x"7f", -- $058a7
          22696 => x"7f", -- $058a8
          22697 => x"7f", -- $058a9
          22698 => x"7f", -- $058aa
          22699 => x"7f", -- $058ab
          22700 => x"7f", -- $058ac
          22701 => x"7f", -- $058ad
          22702 => x"7f", -- $058ae
          22703 => x"7f", -- $058af
          22704 => x"7f", -- $058b0
          22705 => x"7f", -- $058b1
          22706 => x"7f", -- $058b2
          22707 => x"7f", -- $058b3
          22708 => x"7f", -- $058b4
          22709 => x"7f", -- $058b5
          22710 => x"7f", -- $058b6
          22711 => x"7f", -- $058b7
          22712 => x"7e", -- $058b8
          22713 => x"7e", -- $058b9
          22714 => x"7f", -- $058ba
          22715 => x"7f", -- $058bb
          22716 => x"7e", -- $058bc
          22717 => x"7f", -- $058bd
          22718 => x"7f", -- $058be
          22719 => x"7f", -- $058bf
          22720 => x"7e", -- $058c0
          22721 => x"7e", -- $058c1
          22722 => x"7e", -- $058c2
          22723 => x"7e", -- $058c3
          22724 => x"7e", -- $058c4
          22725 => x"7e", -- $058c5
          22726 => x"7e", -- $058c6
          22727 => x"7f", -- $058c7
          22728 => x"7f", -- $058c8
          22729 => x"7f", -- $058c9
          22730 => x"7f", -- $058ca
          22731 => x"7e", -- $058cb
          22732 => x"7e", -- $058cc
          22733 => x"7e", -- $058cd
          22734 => x"7e", -- $058ce
          22735 => x"7e", -- $058cf
          22736 => x"7e", -- $058d0
          22737 => x"7e", -- $058d1
          22738 => x"7e", -- $058d2
          22739 => x"7e", -- $058d3
          22740 => x"7e", -- $058d4
          22741 => x"7e", -- $058d5
          22742 => x"7e", -- $058d6
          22743 => x"7e", -- $058d7
          22744 => x"7e", -- $058d8
          22745 => x"7e", -- $058d9
          22746 => x"7e", -- $058da
          22747 => x"7e", -- $058db
          22748 => x"7e", -- $058dc
          22749 => x"7e", -- $058dd
          22750 => x"7e", -- $058de
          22751 => x"7e", -- $058df
          22752 => x"7e", -- $058e0
          22753 => x"7e", -- $058e1
          22754 => x"7e", -- $058e2
          22755 => x"7f", -- $058e3
          22756 => x"7f", -- $058e4
          22757 => x"7e", -- $058e5
          22758 => x"7f", -- $058e6
          22759 => x"7e", -- $058e7
          22760 => x"7e", -- $058e8
          22761 => x"7e", -- $058e9
          22762 => x"7e", -- $058ea
          22763 => x"7e", -- $058eb
          22764 => x"7e", -- $058ec
          22765 => x"7e", -- $058ed
          22766 => x"7e", -- $058ee
          22767 => x"7e", -- $058ef
          22768 => x"7e", -- $058f0
          22769 => x"7e", -- $058f1
          22770 => x"7e", -- $058f2
          22771 => x"7e", -- $058f3
          22772 => x"7e", -- $058f4
          22773 => x"7e", -- $058f5
          22774 => x"7e", -- $058f6
          22775 => x"7e", -- $058f7
          22776 => x"7e", -- $058f8
          22777 => x"7e", -- $058f9
          22778 => x"7f", -- $058fa
          22779 => x"7f", -- $058fb
          22780 => x"7f", -- $058fc
          22781 => x"7f", -- $058fd
          22782 => x"7f", -- $058fe
          22783 => x"7f", -- $058ff
          22784 => x"7f", -- $05900
          22785 => x"7f", -- $05901
          22786 => x"7f", -- $05902
          22787 => x"7f", -- $05903
          22788 => x"7f", -- $05904
          22789 => x"7f", -- $05905
          22790 => x"7f", -- $05906
          22791 => x"7f", -- $05907
          22792 => x"7f", -- $05908
          22793 => x"7f", -- $05909
          22794 => x"7f", -- $0590a
          22795 => x"7f", -- $0590b
          22796 => x"7f", -- $0590c
          22797 => x"7f", -- $0590d
          22798 => x"7f", -- $0590e
          22799 => x"7f", -- $0590f
          22800 => x"7f", -- $05910
          22801 => x"7f", -- $05911
          22802 => x"7f", -- $05912
          22803 => x"7f", -- $05913
          22804 => x"7f", -- $05914
          22805 => x"80", -- $05915
          22806 => x"80", -- $05916
          22807 => x"80", -- $05917
          22808 => x"80", -- $05918
          22809 => x"80", -- $05919
          22810 => x"80", -- $0591a
          22811 => x"80", -- $0591b
          22812 => x"80", -- $0591c
          22813 => x"80", -- $0591d
          22814 => x"80", -- $0591e
          22815 => x"80", -- $0591f
          22816 => x"80", -- $05920
          22817 => x"80", -- $05921
          22818 => x"80", -- $05922
          22819 => x"80", -- $05923
          22820 => x"80", -- $05924
          22821 => x"80", -- $05925
          22822 => x"80", -- $05926
          22823 => x"80", -- $05927
          22824 => x"80", -- $05928
          22825 => x"80", -- $05929
          22826 => x"80", -- $0592a
          22827 => x"80", -- $0592b
          22828 => x"80", -- $0592c
          22829 => x"80", -- $0592d
          22830 => x"80", -- $0592e
          22831 => x"80", -- $0592f
          22832 => x"80", -- $05930
          22833 => x"80", -- $05931
          22834 => x"80", -- $05932
          22835 => x"80", -- $05933
          22836 => x"80", -- $05934
          22837 => x"80", -- $05935
          22838 => x"80", -- $05936
          22839 => x"80", -- $05937
          22840 => x"80", -- $05938
          22841 => x"80", -- $05939
          22842 => x"80", -- $0593a
          22843 => x"80", -- $0593b
          22844 => x"80", -- $0593c
          22845 => x"80", -- $0593d
          22846 => x"80", -- $0593e
          22847 => x"80", -- $0593f
          22848 => x"80", -- $05940
          22849 => x"80", -- $05941
          22850 => x"80", -- $05942
          22851 => x"80", -- $05943
          22852 => x"80", -- $05944
          22853 => x"80", -- $05945
          22854 => x"80", -- $05946
          22855 => x"80", -- $05947
          22856 => x"80", -- $05948
          22857 => x"80", -- $05949
          22858 => x"80", -- $0594a
          22859 => x"80", -- $0594b
          22860 => x"80", -- $0594c
          22861 => x"80", -- $0594d
          22862 => x"80", -- $0594e
          22863 => x"80", -- $0594f
          22864 => x"80", -- $05950
          22865 => x"80", -- $05951
          22866 => x"80", -- $05952
          22867 => x"80", -- $05953
          22868 => x"80", -- $05954
          22869 => x"80", -- $05955
          22870 => x"80", -- $05956
          22871 => x"80", -- $05957
          22872 => x"80", -- $05958
          22873 => x"80", -- $05959
          22874 => x"80", -- $0595a
          22875 => x"80", -- $0595b
          22876 => x"80", -- $0595c
          22877 => x"80", -- $0595d
          22878 => x"80", -- $0595e
          22879 => x"80", -- $0595f
          22880 => x"80", -- $05960
          22881 => x"80", -- $05961
          22882 => x"80", -- $05962
          22883 => x"80", -- $05963
          22884 => x"80", -- $05964
          22885 => x"80", -- $05965
          22886 => x"80", -- $05966
          22887 => x"80", -- $05967
          22888 => x"80", -- $05968
          22889 => x"80", -- $05969
          22890 => x"80", -- $0596a
          22891 => x"80", -- $0596b
          22892 => x"80", -- $0596c
          22893 => x"80", -- $0596d
          22894 => x"80", -- $0596e
          22895 => x"80", -- $0596f
          22896 => x"80", -- $05970
          22897 => x"80", -- $05971
          22898 => x"80", -- $05972
          22899 => x"80", -- $05973
          22900 => x"80", -- $05974
          22901 => x"80", -- $05975
          22902 => x"80", -- $05976
          22903 => x"80", -- $05977
          22904 => x"80", -- $05978
          22905 => x"80", -- $05979
          22906 => x"80", -- $0597a
          22907 => x"80", -- $0597b
          22908 => x"80", -- $0597c
          22909 => x"80", -- $0597d
          22910 => x"80", -- $0597e
          22911 => x"80", -- $0597f
          22912 => x"80", -- $05980
          22913 => x"80", -- $05981
          22914 => x"80", -- $05982
          22915 => x"80", -- $05983
          22916 => x"80", -- $05984
          22917 => x"80", -- $05985
          22918 => x"80", -- $05986
          22919 => x"80", -- $05987
          22920 => x"80", -- $05988
          22921 => x"80", -- $05989
          22922 => x"80", -- $0598a
          22923 => x"80", -- $0598b
          22924 => x"80", -- $0598c
          22925 => x"80", -- $0598d
          22926 => x"80", -- $0598e
          22927 => x"80", -- $0598f
          22928 => x"80", -- $05990
          22929 => x"80", -- $05991
          22930 => x"80", -- $05992
          22931 => x"80", -- $05993
          22932 => x"80", -- $05994
          22933 => x"80", -- $05995
          22934 => x"80", -- $05996
          22935 => x"80", -- $05997
          22936 => x"80", -- $05998
          22937 => x"80", -- $05999
          22938 => x"80", -- $0599a
          22939 => x"80", -- $0599b
          22940 => x"80", -- $0599c
          22941 => x"80", -- $0599d
          22942 => x"80", -- $0599e
          22943 => x"80", -- $0599f
          22944 => x"80", -- $059a0
          22945 => x"80", -- $059a1
          22946 => x"80", -- $059a2
          22947 => x"80", -- $059a3
          22948 => x"80", -- $059a4
          22949 => x"80", -- $059a5
          22950 => x"80", -- $059a6
          22951 => x"80", -- $059a7
          22952 => x"80", -- $059a8
          22953 => x"80", -- $059a9
          22954 => x"80", -- $059aa
          22955 => x"80", -- $059ab
          22956 => x"80", -- $059ac
          22957 => x"80", -- $059ad
          22958 => x"80", -- $059ae
          22959 => x"80", -- $059af
          22960 => x"80", -- $059b0
          22961 => x"80", -- $059b1
          22962 => x"80", -- $059b2
          22963 => x"80", -- $059b3
          22964 => x"80", -- $059b4
          22965 => x"80", -- $059b5
          22966 => x"80", -- $059b6
          22967 => x"80", -- $059b7
          22968 => x"80", -- $059b8
          22969 => x"80", -- $059b9
          22970 => x"80", -- $059ba
          22971 => x"80", -- $059bb
          22972 => x"80", -- $059bc
          22973 => x"80", -- $059bd
          22974 => x"80", -- $059be
          22975 => x"80", -- $059bf
          22976 => x"80", -- $059c0
          22977 => x"80", -- $059c1
          22978 => x"80", -- $059c2
          22979 => x"80", -- $059c3
          22980 => x"80", -- $059c4
          22981 => x"80", -- $059c5
          22982 => x"80", -- $059c6
          22983 => x"80", -- $059c7
          22984 => x"80", -- $059c8
          22985 => x"80", -- $059c9
          22986 => x"80", -- $059ca
          22987 => x"80", -- $059cb
          22988 => x"80", -- $059cc
          22989 => x"80", -- $059cd
          22990 => x"80", -- $059ce
          22991 => x"80", -- $059cf
          22992 => x"80", -- $059d0
          22993 => x"80", -- $059d1
          22994 => x"80", -- $059d2
          22995 => x"80", -- $059d3
          22996 => x"80", -- $059d4
          22997 => x"80", -- $059d5
          22998 => x"80", -- $059d6
          22999 => x"80", -- $059d7
          23000 => x"80", -- $059d8
          23001 => x"80", -- $059d9
          23002 => x"80", -- $059da
          23003 => x"80", -- $059db
          23004 => x"80", -- $059dc
          23005 => x"80", -- $059dd
          23006 => x"80", -- $059de
          23007 => x"80", -- $059df
          23008 => x"80", -- $059e0
          23009 => x"80", -- $059e1
          23010 => x"80", -- $059e2
          23011 => x"80", -- $059e3
          23012 => x"80", -- $059e4
          23013 => x"80", -- $059e5
          23014 => x"80", -- $059e6
          23015 => x"80", -- $059e7
          23016 => x"80", -- $059e8
          23017 => x"80", -- $059e9
          23018 => x"81", -- $059ea
          23019 => x"81", -- $059eb
          23020 => x"81", -- $059ec
          23021 => x"81", -- $059ed
          23022 => x"81", -- $059ee
          23023 => x"81", -- $059ef
          23024 => x"81", -- $059f0
          23025 => x"81", -- $059f1
          23026 => x"81", -- $059f2
          23027 => x"81", -- $059f3
          23028 => x"81", -- $059f4
          23029 => x"81", -- $059f5
          23030 => x"81", -- $059f6
          23031 => x"81", -- $059f7
          23032 => x"81", -- $059f8
          23033 => x"81", -- $059f9
          23034 => x"81", -- $059fa
          23035 => x"81", -- $059fb
          23036 => x"81", -- $059fc
          23037 => x"81", -- $059fd
          23038 => x"81", -- $059fe
          23039 => x"81", -- $059ff
          23040 => x"81", -- $05a00
          23041 => x"81", -- $05a01
          23042 => x"81", -- $05a02
          23043 => x"81", -- $05a03
          23044 => x"81", -- $05a04
          23045 => x"81", -- $05a05
          23046 => x"81", -- $05a06
          23047 => x"81", -- $05a07
          23048 => x"81", -- $05a08
          23049 => x"81", -- $05a09
          23050 => x"81", -- $05a0a
          23051 => x"81", -- $05a0b
          23052 => x"81", -- $05a0c
          23053 => x"81", -- $05a0d
          23054 => x"81", -- $05a0e
          23055 => x"81", -- $05a0f
          23056 => x"81", -- $05a10
          23057 => x"81", -- $05a11
          23058 => x"81", -- $05a12
          23059 => x"81", -- $05a13
          23060 => x"81", -- $05a14
          23061 => x"81", -- $05a15
          23062 => x"81", -- $05a16
          23063 => x"81", -- $05a17
          23064 => x"81", -- $05a18
          23065 => x"81", -- $05a19
          23066 => x"81", -- $05a1a
          23067 => x"81", -- $05a1b
          23068 => x"81", -- $05a1c
          23069 => x"81", -- $05a1d
          23070 => x"81", -- $05a1e
          23071 => x"81", -- $05a1f
          23072 => x"81", -- $05a20
          23073 => x"81", -- $05a21
          23074 => x"81", -- $05a22
          23075 => x"81", -- $05a23
          23076 => x"81", -- $05a24
          23077 => x"81", -- $05a25
          23078 => x"81", -- $05a26
          23079 => x"81", -- $05a27
          23080 => x"81", -- $05a28
          23081 => x"81", -- $05a29
          23082 => x"81", -- $05a2a
          23083 => x"81", -- $05a2b
          23084 => x"81", -- $05a2c
          23085 => x"81", -- $05a2d
          23086 => x"81", -- $05a2e
          23087 => x"81", -- $05a2f
          23088 => x"81", -- $05a30
          23089 => x"81", -- $05a31
          23090 => x"81", -- $05a32
          23091 => x"81", -- $05a33
          23092 => x"81", -- $05a34
          23093 => x"81", -- $05a35
          23094 => x"81", -- $05a36
          23095 => x"81", -- $05a37
          23096 => x"81", -- $05a38
          23097 => x"81", -- $05a39
          23098 => x"81", -- $05a3a
          23099 => x"81", -- $05a3b
          23100 => x"81", -- $05a3c
          23101 => x"81", -- $05a3d
          23102 => x"81", -- $05a3e
          23103 => x"81", -- $05a3f
          23104 => x"81", -- $05a40
          23105 => x"81", -- $05a41
          23106 => x"81", -- $05a42
          23107 => x"81", -- $05a43
          23108 => x"81", -- $05a44
          23109 => x"81", -- $05a45
          23110 => x"81", -- $05a46
          23111 => x"81", -- $05a47
          23112 => x"80", -- $05a48
          23113 => x"80", -- $05a49
          23114 => x"81", -- $05a4a
          23115 => x"81", -- $05a4b
          23116 => x"81", -- $05a4c
          23117 => x"81", -- $05a4d
          23118 => x"81", -- $05a4e
          23119 => x"81", -- $05a4f
          23120 => x"81", -- $05a50
          23121 => x"81", -- $05a51
          23122 => x"81", -- $05a52
          23123 => x"81", -- $05a53
          23124 => x"81", -- $05a54
          23125 => x"81", -- $05a55
          23126 => x"81", -- $05a56
          23127 => x"81", -- $05a57
          23128 => x"81", -- $05a58
          23129 => x"81", -- $05a59
          23130 => x"81", -- $05a5a
          23131 => x"81", -- $05a5b
          23132 => x"81", -- $05a5c
          23133 => x"81", -- $05a5d
          23134 => x"81", -- $05a5e
          23135 => x"81", -- $05a5f
          23136 => x"81", -- $05a60
          23137 => x"81", -- $05a61
          23138 => x"81", -- $05a62
          23139 => x"81", -- $05a63
          23140 => x"80", -- $05a64
          23141 => x"81", -- $05a65
          23142 => x"81", -- $05a66
          23143 => x"81", -- $05a67
          23144 => x"81", -- $05a68
          23145 => x"81", -- $05a69
          23146 => x"81", -- $05a6a
          23147 => x"81", -- $05a6b
          23148 => x"81", -- $05a6c
          23149 => x"81", -- $05a6d
          23150 => x"81", -- $05a6e
          23151 => x"81", -- $05a6f
          23152 => x"81", -- $05a70
          23153 => x"81", -- $05a71
          23154 => x"81", -- $05a72
          23155 => x"81", -- $05a73
          23156 => x"81", -- $05a74
          23157 => x"80", -- $05a75
          23158 => x"81", -- $05a76
          23159 => x"81", -- $05a77
          23160 => x"81", -- $05a78
          23161 => x"81", -- $05a79
          23162 => x"81", -- $05a7a
          23163 => x"81", -- $05a7b
          23164 => x"81", -- $05a7c
          23165 => x"80", -- $05a7d
          23166 => x"80", -- $05a7e
          23167 => x"81", -- $05a7f
          23168 => x"81", -- $05a80
          23169 => x"81", -- $05a81
          23170 => x"81", -- $05a82
          23171 => x"81", -- $05a83
          23172 => x"81", -- $05a84
          23173 => x"81", -- $05a85
          23174 => x"81", -- $05a86
          23175 => x"81", -- $05a87
          23176 => x"81", -- $05a88
          23177 => x"81", -- $05a89
          23178 => x"81", -- $05a8a
          23179 => x"81", -- $05a8b
          23180 => x"81", -- $05a8c
          23181 => x"81", -- $05a8d
          23182 => x"81", -- $05a8e
          23183 => x"81", -- $05a8f
          23184 => x"81", -- $05a90
          23185 => x"81", -- $05a91
          23186 => x"81", -- $05a92
          23187 => x"81", -- $05a93
          23188 => x"81", -- $05a94
          23189 => x"81", -- $05a95
          23190 => x"81", -- $05a96
          23191 => x"81", -- $05a97
          23192 => x"81", -- $05a98
          23193 => x"81", -- $05a99
          23194 => x"81", -- $05a9a
          23195 => x"81", -- $05a9b
          23196 => x"81", -- $05a9c
          23197 => x"81", -- $05a9d
          23198 => x"81", -- $05a9e
          23199 => x"81", -- $05a9f
          23200 => x"81", -- $05aa0
          23201 => x"81", -- $05aa1
          23202 => x"81", -- $05aa2
          23203 => x"81", -- $05aa3
          23204 => x"81", -- $05aa4
          23205 => x"81", -- $05aa5
          23206 => x"81", -- $05aa6
          23207 => x"81", -- $05aa7
          23208 => x"81", -- $05aa8
          23209 => x"81", -- $05aa9
          23210 => x"81", -- $05aaa
          23211 => x"81", -- $05aab
          23212 => x"81", -- $05aac
          23213 => x"81", -- $05aad
          23214 => x"81", -- $05aae
          23215 => x"81", -- $05aaf
          23216 => x"81", -- $05ab0
          23217 => x"81", -- $05ab1
          23218 => x"81", -- $05ab2
          23219 => x"81", -- $05ab3
          23220 => x"81", -- $05ab4
          23221 => x"81", -- $05ab5
          23222 => x"81", -- $05ab6
          23223 => x"81", -- $05ab7
          23224 => x"81", -- $05ab8
          23225 => x"81", -- $05ab9
          23226 => x"81", -- $05aba
          23227 => x"81", -- $05abb
          23228 => x"81", -- $05abc
          23229 => x"81", -- $05abd
          23230 => x"81", -- $05abe
          23231 => x"81", -- $05abf
          23232 => x"81", -- $05ac0
          23233 => x"81", -- $05ac1
          23234 => x"81", -- $05ac2
          23235 => x"81", -- $05ac3
          23236 => x"81", -- $05ac4
          23237 => x"81", -- $05ac5
          23238 => x"81", -- $05ac6
          23239 => x"81", -- $05ac7
          23240 => x"81", -- $05ac8
          23241 => x"81", -- $05ac9
          23242 => x"81", -- $05aca
          23243 => x"81", -- $05acb
          23244 => x"80", -- $05acc
          23245 => x"80", -- $05acd
          23246 => x"80", -- $05ace
          23247 => x"80", -- $05acf
          23248 => x"80", -- $05ad0
          23249 => x"80", -- $05ad1
          23250 => x"80", -- $05ad2
          23251 => x"81", -- $05ad3
          23252 => x"80", -- $05ad4
          23253 => x"80", -- $05ad5
          23254 => x"80", -- $05ad6
          23255 => x"80", -- $05ad7
          23256 => x"80", -- $05ad8
          23257 => x"80", -- $05ad9
          23258 => x"80", -- $05ada
          23259 => x"80", -- $05adb
          23260 => x"80", -- $05adc
          23261 => x"80", -- $05add
          23262 => x"80", -- $05ade
          23263 => x"80", -- $05adf
          23264 => x"80", -- $05ae0
          23265 => x"80", -- $05ae1
          23266 => x"80", -- $05ae2
          23267 => x"80", -- $05ae3
          23268 => x"80", -- $05ae4
          23269 => x"80", -- $05ae5
          23270 => x"80", -- $05ae6
          23271 => x"80", -- $05ae7
          23272 => x"80", -- $05ae8
          23273 => x"80", -- $05ae9
          23274 => x"80", -- $05aea
          23275 => x"80", -- $05aeb
          23276 => x"80", -- $05aec
          23277 => x"80", -- $05aed
          23278 => x"80", -- $05aee
          23279 => x"80", -- $05aef
          23280 => x"80", -- $05af0
          23281 => x"80", -- $05af1
          23282 => x"80", -- $05af2
          23283 => x"80", -- $05af3
          23284 => x"80", -- $05af4
          23285 => x"80", -- $05af5
          23286 => x"80", -- $05af6
          23287 => x"80", -- $05af7
          23288 => x"80", -- $05af8
          23289 => x"80", -- $05af9
          23290 => x"80", -- $05afa
          23291 => x"80", -- $05afb
          23292 => x"80", -- $05afc
          23293 => x"80", -- $05afd
          23294 => x"80", -- $05afe
          23295 => x"80", -- $05aff
          23296 => x"80", -- $05b00
          23297 => x"80", -- $05b01
          23298 => x"80", -- $05b02
          23299 => x"80", -- $05b03
          23300 => x"80", -- $05b04
          23301 => x"80", -- $05b05
          23302 => x"80", -- $05b06
          23303 => x"80", -- $05b07
          23304 => x"80", -- $05b08
          23305 => x"80", -- $05b09
          23306 => x"80", -- $05b0a
          23307 => x"80", -- $05b0b
          23308 => x"80", -- $05b0c
          23309 => x"80", -- $05b0d
          23310 => x"80", -- $05b0e
          23311 => x"80", -- $05b0f
          23312 => x"80", -- $05b10
          23313 => x"80", -- $05b11
          23314 => x"80", -- $05b12
          23315 => x"80", -- $05b13
          23316 => x"80", -- $05b14
          23317 => x"80", -- $05b15
          23318 => x"80", -- $05b16
          23319 => x"80", -- $05b17
          23320 => x"80", -- $05b18
          23321 => x"80", -- $05b19
          23322 => x"80", -- $05b1a
          23323 => x"80", -- $05b1b
          23324 => x"80", -- $05b1c
          23325 => x"80", -- $05b1d
          23326 => x"80", -- $05b1e
          23327 => x"80", -- $05b1f
          23328 => x"80", -- $05b20
          23329 => x"80", -- $05b21
          23330 => x"80", -- $05b22
          23331 => x"80", -- $05b23
          23332 => x"80", -- $05b24
          23333 => x"80", -- $05b25
          23334 => x"80", -- $05b26
          23335 => x"80", -- $05b27
          23336 => x"80", -- $05b28
          23337 => x"80", -- $05b29
          23338 => x"80", -- $05b2a
          23339 => x"80", -- $05b2b
          23340 => x"80", -- $05b2c
          23341 => x"80", -- $05b2d
          23342 => x"80", -- $05b2e
          23343 => x"80", -- $05b2f
          23344 => x"80", -- $05b30
          23345 => x"80", -- $05b31
          23346 => x"80", -- $05b32
          23347 => x"80", -- $05b33
          23348 => x"80", -- $05b34
          23349 => x"80", -- $05b35
          23350 => x"80", -- $05b36
          23351 => x"80", -- $05b37
          23352 => x"80", -- $05b38
          23353 => x"80", -- $05b39
          23354 => x"80", -- $05b3a
          23355 => x"80", -- $05b3b
          23356 => x"80", -- $05b3c
          23357 => x"80", -- $05b3d
          23358 => x"80", -- $05b3e
          23359 => x"80", -- $05b3f
          23360 => x"80", -- $05b40
          23361 => x"7f", -- $05b41
          23362 => x"7f", -- $05b42
          23363 => x"7f", -- $05b43
          23364 => x"7f", -- $05b44
          23365 => x"7f", -- $05b45
          23366 => x"7f", -- $05b46
          23367 => x"7f", -- $05b47
          23368 => x"7f", -- $05b48
          23369 => x"7f", -- $05b49
          23370 => x"7f", -- $05b4a
          23371 => x"7f", -- $05b4b
          23372 => x"7f", -- $05b4c
          23373 => x"7f", -- $05b4d
          23374 => x"7f", -- $05b4e
          23375 => x"7f", -- $05b4f
          23376 => x"7f", -- $05b50
          23377 => x"7f", -- $05b51
          23378 => x"7f", -- $05b52
          23379 => x"7f", -- $05b53
          23380 => x"7f", -- $05b54
          23381 => x"7f", -- $05b55
          23382 => x"7f", -- $05b56
          23383 => x"7f", -- $05b57
          23384 => x"7f", -- $05b58
          23385 => x"7f", -- $05b59
          23386 => x"7f", -- $05b5a
          23387 => x"7f", -- $05b5b
          23388 => x"7f", -- $05b5c
          23389 => x"7f", -- $05b5d
          23390 => x"7f", -- $05b5e
          23391 => x"7f", -- $05b5f
          23392 => x"7f", -- $05b60
          23393 => x"7f", -- $05b61
          23394 => x"7f", -- $05b62
          23395 => x"7f", -- $05b63
          23396 => x"7f", -- $05b64
          23397 => x"7f", -- $05b65
          23398 => x"7f", -- $05b66
          23399 => x"7f", -- $05b67
          23400 => x"7f", -- $05b68
          23401 => x"7f", -- $05b69
          23402 => x"7f", -- $05b6a
          23403 => x"7f", -- $05b6b
          23404 => x"7f", -- $05b6c
          23405 => x"7f", -- $05b6d
          23406 => x"7f", -- $05b6e
          23407 => x"7f", -- $05b6f
          23408 => x"7f", -- $05b70
          23409 => x"7f", -- $05b71
          23410 => x"7f", -- $05b72
          23411 => x"7f", -- $05b73
          23412 => x"7f", -- $05b74
          23413 => x"7f", -- $05b75
          23414 => x"7f", -- $05b76
          23415 => x"7f", -- $05b77
          23416 => x"7f", -- $05b78
          23417 => x"7f", -- $05b79
          23418 => x"7f", -- $05b7a
          23419 => x"7f", -- $05b7b
          23420 => x"7f", -- $05b7c
          23421 => x"7f", -- $05b7d
          23422 => x"7f", -- $05b7e
          23423 => x"7f", -- $05b7f
          23424 => x"7f", -- $05b80
          23425 => x"7f", -- $05b81
          23426 => x"7f", -- $05b82
          23427 => x"7f", -- $05b83
          23428 => x"7f", -- $05b84
          23429 => x"7f", -- $05b85
          23430 => x"7f", -- $05b86
          23431 => x"7f", -- $05b87
          23432 => x"7f", -- $05b88
          23433 => x"7f", -- $05b89
          23434 => x"7f", -- $05b8a
          23435 => x"7f", -- $05b8b
          23436 => x"7f", -- $05b8c
          23437 => x"7f", -- $05b8d
          23438 => x"7f", -- $05b8e
          23439 => x"7f", -- $05b8f
          23440 => x"7f", -- $05b90
          23441 => x"7f", -- $05b91
          23442 => x"7f", -- $05b92
          23443 => x"7f", -- $05b93
          23444 => x"7f", -- $05b94
          23445 => x"7f", -- $05b95
          23446 => x"7f", -- $05b96
          23447 => x"7f", -- $05b97
          23448 => x"80", -- $05b98
          23449 => x"7f", -- $05b99
          23450 => x"7f", -- $05b9a
          23451 => x"7f", -- $05b9b
          23452 => x"7f", -- $05b9c
          23453 => x"7f", -- $05b9d
          23454 => x"7f", -- $05b9e
          23455 => x"7f", -- $05b9f
          23456 => x"7f", -- $05ba0
          23457 => x"7f", -- $05ba1
          23458 => x"7f", -- $05ba2
          23459 => x"7f", -- $05ba3
          23460 => x"7f", -- $05ba4
          23461 => x"80", -- $05ba5
          23462 => x"7f", -- $05ba6
          23463 => x"7f", -- $05ba7
          23464 => x"7f", -- $05ba8
          23465 => x"7f", -- $05ba9
          23466 => x"7f", -- $05baa
          23467 => x"7f", -- $05bab
          23468 => x"7f", -- $05bac
          23469 => x"7f", -- $05bad
          23470 => x"7f", -- $05bae
          23471 => x"7f", -- $05baf
          23472 => x"7f", -- $05bb0
          23473 => x"7f", -- $05bb1
          23474 => x"7f", -- $05bb2
          23475 => x"7f", -- $05bb3
          23476 => x"80", -- $05bb4
          23477 => x"7f", -- $05bb5
          23478 => x"7f", -- $05bb6
          23479 => x"80", -- $05bb7
          23480 => x"80", -- $05bb8
          23481 => x"80", -- $05bb9
          23482 => x"80", -- $05bba
          23483 => x"80", -- $05bbb
          23484 => x"80", -- $05bbc
          23485 => x"80", -- $05bbd
          23486 => x"80", -- $05bbe
          23487 => x"80", -- $05bbf
          23488 => x"80", -- $05bc0
          23489 => x"80", -- $05bc1
          23490 => x"80", -- $05bc2
          23491 => x"80", -- $05bc3
          23492 => x"80", -- $05bc4
          23493 => x"80", -- $05bc5
          23494 => x"80", -- $05bc6
          23495 => x"80", -- $05bc7
          23496 => x"80", -- $05bc8
          23497 => x"80", -- $05bc9
          23498 => x"80", -- $05bca
          23499 => x"80", -- $05bcb
          23500 => x"80", -- $05bcc
          23501 => x"80", -- $05bcd
          23502 => x"80", -- $05bce
          23503 => x"80", -- $05bcf
          23504 => x"80", -- $05bd0
          23505 => x"80", -- $05bd1
          23506 => x"80", -- $05bd2
          23507 => x"80", -- $05bd3
          23508 => x"80", -- $05bd4
          23509 => x"80", -- $05bd5
          23510 => x"80", -- $05bd6
          23511 => x"80", -- $05bd7
          23512 => x"80", -- $05bd8
          23513 => x"80", -- $05bd9
          23514 => x"80", -- $05bda
          23515 => x"80", -- $05bdb
          23516 => x"80", -- $05bdc
          23517 => x"80", -- $05bdd
          23518 => x"80", -- $05bde
          23519 => x"80", -- $05bdf
          23520 => x"7f", -- $05be0
          23521 => x"7f", -- $05be1
          23522 => x"7f", -- $05be2
          23523 => x"7f", -- $05be3
          23524 => x"80", -- $05be4
          23525 => x"80", -- $05be5
          23526 => x"80", -- $05be6
          23527 => x"80", -- $05be7
          23528 => x"80", -- $05be8
          23529 => x"80", -- $05be9
          23530 => x"80", -- $05bea
          23531 => x"80", -- $05beb
          23532 => x"80", -- $05bec
          23533 => x"80", -- $05bed
          23534 => x"80", -- $05bee
          23535 => x"80", -- $05bef
          23536 => x"80", -- $05bf0
          23537 => x"80", -- $05bf1
          23538 => x"80", -- $05bf2
          23539 => x"80", -- $05bf3
          23540 => x"80", -- $05bf4
          23541 => x"80", -- $05bf5
          23542 => x"80", -- $05bf6
          23543 => x"7f", -- $05bf7
          23544 => x"7f", -- $05bf8
          23545 => x"7f", -- $05bf9
          23546 => x"7f", -- $05bfa
          23547 => x"7f", -- $05bfb
          23548 => x"7f", -- $05bfc
          23549 => x"7f", -- $05bfd
          23550 => x"80", -- $05bfe
          23551 => x"80", -- $05bff
          23552 => x"80", -- $05c00
          23553 => x"7f", -- $05c01
          23554 => x"7f", -- $05c02
          23555 => x"7f", -- $05c03
          23556 => x"7f", -- $05c04
          23557 => x"7f", -- $05c05
          23558 => x"7f", -- $05c06
          23559 => x"7f", -- $05c07
          23560 => x"7f", -- $05c08
          23561 => x"7f", -- $05c09
          23562 => x"7f", -- $05c0a
          23563 => x"7f", -- $05c0b
          23564 => x"7f", -- $05c0c
          23565 => x"7f", -- $05c0d
          23566 => x"7f", -- $05c0e
          23567 => x"7f", -- $05c0f
          23568 => x"7f", -- $05c10
          23569 => x"7f", -- $05c11
          23570 => x"7f", -- $05c12
          23571 => x"7f", -- $05c13
          23572 => x"7f", -- $05c14
          23573 => x"7f", -- $05c15
          23574 => x"7f", -- $05c16
          23575 => x"7f", -- $05c17
          23576 => x"7f", -- $05c18
          23577 => x"7f", -- $05c19
          23578 => x"7f", -- $05c1a
          23579 => x"7f", -- $05c1b
          23580 => x"7f", -- $05c1c
          23581 => x"7f", -- $05c1d
          23582 => x"7f", -- $05c1e
          23583 => x"7f", -- $05c1f
          23584 => x"7f", -- $05c20
          23585 => x"7f", -- $05c21
          23586 => x"7f", -- $05c22
          23587 => x"7f", -- $05c23
          23588 => x"7f", -- $05c24
          23589 => x"7f", -- $05c25
          23590 => x"7f", -- $05c26
          23591 => x"7f", -- $05c27
          23592 => x"7f", -- $05c28
          23593 => x"7f", -- $05c29
          23594 => x"7f", -- $05c2a
          23595 => x"7f", -- $05c2b
          23596 => x"7f", -- $05c2c
          23597 => x"7f", -- $05c2d
          23598 => x"7f", -- $05c2e
          23599 => x"7f", -- $05c2f
          23600 => x"7f", -- $05c30
          23601 => x"7f", -- $05c31
          23602 => x"7f", -- $05c32
          23603 => x"7f", -- $05c33
          23604 => x"7f", -- $05c34
          23605 => x"7f", -- $05c35
          23606 => x"7f", -- $05c36
          23607 => x"7f", -- $05c37
          23608 => x"7f", -- $05c38
          23609 => x"7f", -- $05c39
          23610 => x"7f", -- $05c3a
          23611 => x"7f", -- $05c3b
          23612 => x"7f", -- $05c3c
          23613 => x"7f", -- $05c3d
          23614 => x"7f", -- $05c3e
          23615 => x"7f", -- $05c3f
          23616 => x"7f", -- $05c40
          23617 => x"7f", -- $05c41
          23618 => x"7f", -- $05c42
          23619 => x"7f", -- $05c43
          23620 => x"7f", -- $05c44
          23621 => x"7f", -- $05c45
          23622 => x"7f", -- $05c46
          23623 => x"7f", -- $05c47
          23624 => x"7f", -- $05c48
          23625 => x"7f", -- $05c49
          23626 => x"7f", -- $05c4a
          23627 => x"7f", -- $05c4b
          23628 => x"7f", -- $05c4c
          23629 => x"7f", -- $05c4d
          23630 => x"7f", -- $05c4e
          23631 => x"7f", -- $05c4f
          23632 => x"7f", -- $05c50
          23633 => x"7f", -- $05c51
          23634 => x"7f", -- $05c52
          23635 => x"7f", -- $05c53
          23636 => x"7f", -- $05c54
          23637 => x"7f", -- $05c55
          23638 => x"80", -- $05c56
          23639 => x"80", -- $05c57
          23640 => x"80", -- $05c58
          23641 => x"80", -- $05c59
          23642 => x"80", -- $05c5a
          23643 => x"80", -- $05c5b
          23644 => x"80", -- $05c5c
          23645 => x"80", -- $05c5d
          23646 => x"80", -- $05c5e
          23647 => x"80", -- $05c5f
          23648 => x"80", -- $05c60
          23649 => x"80", -- $05c61
          23650 => x"80", -- $05c62
          23651 => x"80", -- $05c63
          23652 => x"80", -- $05c64
          23653 => x"80", -- $05c65
          23654 => x"80", -- $05c66
          23655 => x"80", -- $05c67
          23656 => x"80", -- $05c68
          23657 => x"80", -- $05c69
          23658 => x"80", -- $05c6a
          23659 => x"80", -- $05c6b
          23660 => x"80", -- $05c6c
          23661 => x"80", -- $05c6d
          23662 => x"80", -- $05c6e
          23663 => x"80", -- $05c6f
          23664 => x"80", -- $05c70
          23665 => x"80", -- $05c71
          23666 => x"80", -- $05c72
          23667 => x"80", -- $05c73
          23668 => x"80", -- $05c74
          23669 => x"80", -- $05c75
          23670 => x"80", -- $05c76
          23671 => x"80", -- $05c77
          23672 => x"80", -- $05c78
          23673 => x"80", -- $05c79
          23674 => x"80", -- $05c7a
          23675 => x"80", -- $05c7b
          23676 => x"80", -- $05c7c
          23677 => x"80", -- $05c7d
          23678 => x"80", -- $05c7e
          23679 => x"80", -- $05c7f
          23680 => x"80", -- $05c80
          23681 => x"80", -- $05c81
          23682 => x"80", -- $05c82
          23683 => x"80", -- $05c83
          23684 => x"80", -- $05c84
          23685 => x"80", -- $05c85
          23686 => x"80", -- $05c86
          23687 => x"80", -- $05c87
          23688 => x"80", -- $05c88
          23689 => x"80", -- $05c89
          23690 => x"80", -- $05c8a
          23691 => x"80", -- $05c8b
          23692 => x"80", -- $05c8c
          23693 => x"80", -- $05c8d
          23694 => x"80", -- $05c8e
          23695 => x"80", -- $05c8f
          23696 => x"80", -- $05c90
          23697 => x"80", -- $05c91
          23698 => x"80", -- $05c92
          23699 => x"80", -- $05c93
          23700 => x"80", -- $05c94
          23701 => x"80", -- $05c95
          23702 => x"80", -- $05c96
          23703 => x"80", -- $05c97
          23704 => x"80", -- $05c98
          23705 => x"80", -- $05c99
          23706 => x"80", -- $05c9a
          23707 => x"80", -- $05c9b
          23708 => x"80", -- $05c9c
          23709 => x"80", -- $05c9d
          23710 => x"80", -- $05c9e
          23711 => x"80", -- $05c9f
          23712 => x"80", -- $05ca0
          23713 => x"80", -- $05ca1
          23714 => x"80", -- $05ca2
          23715 => x"80", -- $05ca3
          23716 => x"80", -- $05ca4
          23717 => x"80", -- $05ca5
          23718 => x"80", -- $05ca6
          23719 => x"80", -- $05ca7
          23720 => x"80", -- $05ca8
          23721 => x"80", -- $05ca9
          23722 => x"80", -- $05caa
          23723 => x"80", -- $05cab
          23724 => x"80", -- $05cac
          23725 => x"80", -- $05cad
          23726 => x"80", -- $05cae
          23727 => x"80", -- $05caf
          23728 => x"80", -- $05cb0
          23729 => x"80", -- $05cb1
          23730 => x"80", -- $05cb2
          23731 => x"80", -- $05cb3
          23732 => x"80", -- $05cb4
          23733 => x"80", -- $05cb5
          23734 => x"80", -- $05cb6
          23735 => x"80", -- $05cb7
          23736 => x"80", -- $05cb8
          23737 => x"80", -- $05cb9
          23738 => x"80", -- $05cba
          23739 => x"80", -- $05cbb
          23740 => x"80", -- $05cbc
          23741 => x"80", -- $05cbd
          23742 => x"80", -- $05cbe
          23743 => x"80", -- $05cbf
          23744 => x"80", -- $05cc0
          23745 => x"80", -- $05cc1
          23746 => x"80", -- $05cc2
          23747 => x"80", -- $05cc3
          23748 => x"80", -- $05cc4
          23749 => x"80", -- $05cc5
          23750 => x"80", -- $05cc6
          23751 => x"80", -- $05cc7
          23752 => x"80", -- $05cc8
          23753 => x"80", -- $05cc9
          23754 => x"80", -- $05cca
          23755 => x"80", -- $05ccb
          23756 => x"81", -- $05ccc
          23757 => x"81", -- $05ccd
          23758 => x"80", -- $05cce
          23759 => x"81", -- $05ccf
          23760 => x"81", -- $05cd0
          23761 => x"81", -- $05cd1
          23762 => x"80", -- $05cd2
          23763 => x"80", -- $05cd3
          23764 => x"80", -- $05cd4
          23765 => x"80", -- $05cd5
          23766 => x"80", -- $05cd6
          23767 => x"80", -- $05cd7
          23768 => x"80", -- $05cd8
          23769 => x"80", -- $05cd9
          23770 => x"80", -- $05cda
          23771 => x"81", -- $05cdb
          23772 => x"81", -- $05cdc
          23773 => x"81", -- $05cdd
          23774 => x"81", -- $05cde
          23775 => x"80", -- $05cdf
          23776 => x"81", -- $05ce0
          23777 => x"81", -- $05ce1
          23778 => x"81", -- $05ce2
          23779 => x"80", -- $05ce3
          23780 => x"81", -- $05ce4
          23781 => x"80", -- $05ce5
          23782 => x"81", -- $05ce6
          23783 => x"81", -- $05ce7
          23784 => x"81", -- $05ce8
          23785 => x"81", -- $05ce9
          23786 => x"81", -- $05cea
          23787 => x"81", -- $05ceb
          23788 => x"81", -- $05cec
          23789 => x"81", -- $05ced
          23790 => x"81", -- $05cee
          23791 => x"81", -- $05cef
          23792 => x"81", -- $05cf0
          23793 => x"81", -- $05cf1
          23794 => x"81", -- $05cf2
          23795 => x"81", -- $05cf3
          23796 => x"81", -- $05cf4
          23797 => x"81", -- $05cf5
          23798 => x"81", -- $05cf6
          23799 => x"81", -- $05cf7
          23800 => x"81", -- $05cf8
          23801 => x"81", -- $05cf9
          23802 => x"81", -- $05cfa
          23803 => x"81", -- $05cfb
          23804 => x"80", -- $05cfc
          23805 => x"80", -- $05cfd
          23806 => x"80", -- $05cfe
          23807 => x"81", -- $05cff
          23808 => x"81", -- $05d00
          23809 => x"81", -- $05d01
          23810 => x"81", -- $05d02
          23811 => x"81", -- $05d03
          23812 => x"81", -- $05d04
          23813 => x"81", -- $05d05
          23814 => x"81", -- $05d06
          23815 => x"81", -- $05d07
          23816 => x"81", -- $05d08
          23817 => x"81", -- $05d09
          23818 => x"80", -- $05d0a
          23819 => x"80", -- $05d0b
          23820 => x"80", -- $05d0c
          23821 => x"80", -- $05d0d
          23822 => x"80", -- $05d0e
          23823 => x"81", -- $05d0f
          23824 => x"81", -- $05d10
          23825 => x"81", -- $05d11
          23826 => x"81", -- $05d12
          23827 => x"81", -- $05d13
          23828 => x"81", -- $05d14
          23829 => x"81", -- $05d15
          23830 => x"81", -- $05d16
          23831 => x"81", -- $05d17
          23832 => x"81", -- $05d18
          23833 => x"81", -- $05d19
          23834 => x"81", -- $05d1a
          23835 => x"81", -- $05d1b
          23836 => x"81", -- $05d1c
          23837 => x"81", -- $05d1d
          23838 => x"81", -- $05d1e
          23839 => x"81", -- $05d1f
          23840 => x"81", -- $05d20
          23841 => x"81", -- $05d21
          23842 => x"81", -- $05d22
          23843 => x"81", -- $05d23
          23844 => x"81", -- $05d24
          23845 => x"81", -- $05d25
          23846 => x"81", -- $05d26
          23847 => x"81", -- $05d27
          23848 => x"81", -- $05d28
          23849 => x"81", -- $05d29
          23850 => x"81", -- $05d2a
          23851 => x"81", -- $05d2b
          23852 => x"81", -- $05d2c
          23853 => x"81", -- $05d2d
          23854 => x"81", -- $05d2e
          23855 => x"81", -- $05d2f
          23856 => x"81", -- $05d30
          23857 => x"81", -- $05d31
          23858 => x"81", -- $05d32
          23859 => x"81", -- $05d33
          23860 => x"81", -- $05d34
          23861 => x"81", -- $05d35
          23862 => x"81", -- $05d36
          23863 => x"81", -- $05d37
          23864 => x"81", -- $05d38
          23865 => x"81", -- $05d39
          23866 => x"81", -- $05d3a
          23867 => x"81", -- $05d3b
          23868 => x"81", -- $05d3c
          23869 => x"81", -- $05d3d
          23870 => x"81", -- $05d3e
          23871 => x"81", -- $05d3f
          23872 => x"81", -- $05d40
          23873 => x"81", -- $05d41
          23874 => x"81", -- $05d42
          23875 => x"81", -- $05d43
          23876 => x"81", -- $05d44
          23877 => x"81", -- $05d45
          23878 => x"81", -- $05d46
          23879 => x"81", -- $05d47
          23880 => x"81", -- $05d48
          23881 => x"81", -- $05d49
          23882 => x"81", -- $05d4a
          23883 => x"81", -- $05d4b
          23884 => x"81", -- $05d4c
          23885 => x"81", -- $05d4d
          23886 => x"81", -- $05d4e
          23887 => x"81", -- $05d4f
          23888 => x"81", -- $05d50
          23889 => x"81", -- $05d51
          23890 => x"81", -- $05d52
          23891 => x"81", -- $05d53
          23892 => x"81", -- $05d54
          23893 => x"81", -- $05d55
          23894 => x"81", -- $05d56
          23895 => x"81", -- $05d57
          23896 => x"81", -- $05d58
          23897 => x"81", -- $05d59
          23898 => x"81", -- $05d5a
          23899 => x"81", -- $05d5b
          23900 => x"81", -- $05d5c
          23901 => x"81", -- $05d5d
          23902 => x"81", -- $05d5e
          23903 => x"81", -- $05d5f
          23904 => x"81", -- $05d60
          23905 => x"81", -- $05d61
          23906 => x"81", -- $05d62
          23907 => x"81", -- $05d63
          23908 => x"81", -- $05d64
          23909 => x"81", -- $05d65
          23910 => x"81", -- $05d66
          23911 => x"81", -- $05d67
          23912 => x"81", -- $05d68
          23913 => x"81", -- $05d69
          23914 => x"81", -- $05d6a
          23915 => x"81", -- $05d6b
          23916 => x"81", -- $05d6c
          23917 => x"81", -- $05d6d
          23918 => x"81", -- $05d6e
          23919 => x"81", -- $05d6f
          23920 => x"81", -- $05d70
          23921 => x"81", -- $05d71
          23922 => x"81", -- $05d72
          23923 => x"81", -- $05d73
          23924 => x"81", -- $05d74
          23925 => x"81", -- $05d75
          23926 => x"81", -- $05d76
          23927 => x"81", -- $05d77
          23928 => x"81", -- $05d78
          23929 => x"81", -- $05d79
          23930 => x"81", -- $05d7a
          23931 => x"81", -- $05d7b
          23932 => x"81", -- $05d7c
          23933 => x"81", -- $05d7d
          23934 => x"81", -- $05d7e
          23935 => x"81", -- $05d7f
          23936 => x"81", -- $05d80
          23937 => x"81", -- $05d81
          23938 => x"81", -- $05d82
          23939 => x"81", -- $05d83
          23940 => x"81", -- $05d84
          23941 => x"81", -- $05d85
          23942 => x"81", -- $05d86
          23943 => x"81", -- $05d87
          23944 => x"81", -- $05d88
          23945 => x"81", -- $05d89
          23946 => x"81", -- $05d8a
          23947 => x"81", -- $05d8b
          23948 => x"80", -- $05d8c
          23949 => x"80", -- $05d8d
          23950 => x"81", -- $05d8e
          23951 => x"80", -- $05d8f
          23952 => x"80", -- $05d90
          23953 => x"80", -- $05d91
          23954 => x"81", -- $05d92
          23955 => x"80", -- $05d93
          23956 => x"80", -- $05d94
          23957 => x"80", -- $05d95
          23958 => x"80", -- $05d96
          23959 => x"80", -- $05d97
          23960 => x"80", -- $05d98
          23961 => x"80", -- $05d99
          23962 => x"80", -- $05d9a
          23963 => x"80", -- $05d9b
          23964 => x"80", -- $05d9c
          23965 => x"80", -- $05d9d
          23966 => x"80", -- $05d9e
          23967 => x"80", -- $05d9f
          23968 => x"80", -- $05da0
          23969 => x"80", -- $05da1
          23970 => x"80", -- $05da2
          23971 => x"80", -- $05da3
          23972 => x"80", -- $05da4
          23973 => x"80", -- $05da5
          23974 => x"80", -- $05da6
          23975 => x"80", -- $05da7
          23976 => x"80", -- $05da8
          23977 => x"80", -- $05da9
          23978 => x"80", -- $05daa
          23979 => x"80", -- $05dab
          23980 => x"80", -- $05dac
          23981 => x"80", -- $05dad
          23982 => x"80", -- $05dae
          23983 => x"80", -- $05daf
          23984 => x"80", -- $05db0
          23985 => x"80", -- $05db1
          23986 => x"80", -- $05db2
          23987 => x"80", -- $05db3
          23988 => x"80", -- $05db4
          23989 => x"80", -- $05db5
          23990 => x"80", -- $05db6
          23991 => x"80", -- $05db7
          23992 => x"80", -- $05db8
          23993 => x"80", -- $05db9
          23994 => x"80", -- $05dba
          23995 => x"80", -- $05dbb
          23996 => x"80", -- $05dbc
          23997 => x"80", -- $05dbd
          23998 => x"80", -- $05dbe
          23999 => x"80", -- $05dbf
          24000 => x"80", -- $05dc0
          24001 => x"80", -- $05dc1
          24002 => x"80", -- $05dc2
          24003 => x"80", -- $05dc3
          24004 => x"80", -- $05dc4
          24005 => x"80", -- $05dc5
          24006 => x"80", -- $05dc6
          24007 => x"80", -- $05dc7
          24008 => x"80", -- $05dc8
          24009 => x"80", -- $05dc9
          24010 => x"80", -- $05dca
          24011 => x"80", -- $05dcb
          24012 => x"80", -- $05dcc
          24013 => x"80", -- $05dcd
          24014 => x"80", -- $05dce
          24015 => x"80", -- $05dcf
          24016 => x"80", -- $05dd0
          24017 => x"80", -- $05dd1
          24018 => x"80", -- $05dd2
          24019 => x"80", -- $05dd3
          24020 => x"80", -- $05dd4
          24021 => x"80", -- $05dd5
          24022 => x"80", -- $05dd6
          24023 => x"80", -- $05dd7
          24024 => x"80", -- $05dd8
          24025 => x"80", -- $05dd9
          24026 => x"80", -- $05dda
          24027 => x"80", -- $05ddb
          24028 => x"80", -- $05ddc
          24029 => x"80", -- $05ddd
          24030 => x"80", -- $05dde
          24031 => x"80", -- $05ddf
          24032 => x"80", -- $05de0
          24033 => x"80", -- $05de1
          24034 => x"80", -- $05de2
          24035 => x"80", -- $05de3
          24036 => x"80", -- $05de4
          24037 => x"80", -- $05de5
          24038 => x"80", -- $05de6
          24039 => x"80", -- $05de7
          24040 => x"80", -- $05de8
          24041 => x"80", -- $05de9
          24042 => x"80", -- $05dea
          24043 => x"80", -- $05deb
          24044 => x"80", -- $05dec
          24045 => x"80", -- $05ded
          24046 => x"80", -- $05dee
          24047 => x"80", -- $05def
          24048 => x"80", -- $05df0
          24049 => x"80", -- $05df1
          24050 => x"80", -- $05df2
          24051 => x"80", -- $05df3
          24052 => x"80", -- $05df4
          24053 => x"80", -- $05df5
          24054 => x"80", -- $05df6
          24055 => x"80", -- $05df7
          24056 => x"80", -- $05df8
          24057 => x"80", -- $05df9
          24058 => x"80", -- $05dfa
          24059 => x"80", -- $05dfb
          24060 => x"80", -- $05dfc
          24061 => x"80", -- $05dfd
          24062 => x"80", -- $05dfe
          24063 => x"80", -- $05dff
          24064 => x"80", -- $05e00
          24065 => x"80", -- $05e01
          24066 => x"80", -- $05e02
          24067 => x"80", -- $05e03
          24068 => x"80", -- $05e04
          24069 => x"80", -- $05e05
          24070 => x"80", -- $05e06
          24071 => x"80", -- $05e07
          24072 => x"80", -- $05e08
          24073 => x"80", -- $05e09
          24074 => x"80", -- $05e0a
          24075 => x"80", -- $05e0b
          24076 => x"80", -- $05e0c
          24077 => x"80", -- $05e0d
          24078 => x"80", -- $05e0e
          24079 => x"80", -- $05e0f
          24080 => x"80", -- $05e10
          24081 => x"80", -- $05e11
          24082 => x"80", -- $05e12
          24083 => x"80", -- $05e13
          24084 => x"80", -- $05e14
          24085 => x"80", -- $05e15
          24086 => x"80", -- $05e16
          24087 => x"80", -- $05e17
          24088 => x"80", -- $05e18
          24089 => x"80", -- $05e19
          24090 => x"80", -- $05e1a
          24091 => x"80", -- $05e1b
          24092 => x"80", -- $05e1c
          24093 => x"80", -- $05e1d
          24094 => x"80", -- $05e1e
          24095 => x"80", -- $05e1f
          24096 => x"80", -- $05e20
          24097 => x"80", -- $05e21
          24098 => x"80", -- $05e22
          24099 => x"80", -- $05e23
          24100 => x"80", -- $05e24
          24101 => x"80", -- $05e25
          24102 => x"80", -- $05e26
          24103 => x"80", -- $05e27
          24104 => x"80", -- $05e28
          24105 => x"80", -- $05e29
          24106 => x"80", -- $05e2a
          24107 => x"80", -- $05e2b
          24108 => x"80", -- $05e2c
          24109 => x"80", -- $05e2d
          24110 => x"80", -- $05e2e
          24111 => x"80", -- $05e2f
          24112 => x"80", -- $05e30
          24113 => x"80", -- $05e31
          24114 => x"80", -- $05e32
          24115 => x"80", -- $05e33
          24116 => x"80", -- $05e34
          24117 => x"80", -- $05e35
          24118 => x"80", -- $05e36
          24119 => x"80", -- $05e37
          24120 => x"80", -- $05e38
          24121 => x"80", -- $05e39
          24122 => x"80", -- $05e3a
          24123 => x"80", -- $05e3b
          24124 => x"80", -- $05e3c
          24125 => x"80", -- $05e3d
          24126 => x"80", -- $05e3e
          24127 => x"80", -- $05e3f
          24128 => x"80", -- $05e40
          24129 => x"80", -- $05e41
          24130 => x"80", -- $05e42
          24131 => x"80", -- $05e43
          24132 => x"80", -- $05e44
          24133 => x"80", -- $05e45
          24134 => x"80", -- $05e46
          24135 => x"80", -- $05e47
          24136 => x"80", -- $05e48
          24137 => x"80", -- $05e49
          24138 => x"80", -- $05e4a
          24139 => x"80", -- $05e4b
          24140 => x"80", -- $05e4c
          24141 => x"80", -- $05e4d
          24142 => x"80", -- $05e4e
          24143 => x"80", -- $05e4f
          24144 => x"80", -- $05e50
          24145 => x"80", -- $05e51
          24146 => x"80", -- $05e52
          24147 => x"80", -- $05e53
          24148 => x"80", -- $05e54
          24149 => x"80", -- $05e55
          24150 => x"80", -- $05e56
          24151 => x"80", -- $05e57
          24152 => x"80", -- $05e58
          24153 => x"80", -- $05e59
          24154 => x"80", -- $05e5a
          24155 => x"80", -- $05e5b
          24156 => x"80", -- $05e5c
          24157 => x"80", -- $05e5d
          24158 => x"80", -- $05e5e
          24159 => x"80", -- $05e5f
          24160 => x"80", -- $05e60
          24161 => x"80", -- $05e61
          24162 => x"80", -- $05e62
          24163 => x"80", -- $05e63
          24164 => x"80", -- $05e64
          24165 => x"80", -- $05e65
          24166 => x"80", -- $05e66
          24167 => x"80", -- $05e67
          24168 => x"80", -- $05e68
          24169 => x"80", -- $05e69
          24170 => x"80", -- $05e6a
          24171 => x"80", -- $05e6b
          24172 => x"80", -- $05e6c
          24173 => x"80", -- $05e6d
          24174 => x"80", -- $05e6e
          24175 => x"80", -- $05e6f
          24176 => x"80", -- $05e70
          24177 => x"80", -- $05e71
          24178 => x"80", -- $05e72
          24179 => x"80", -- $05e73
          24180 => x"80", -- $05e74
          24181 => x"80", -- $05e75
          24182 => x"80", -- $05e76
          24183 => x"80", -- $05e77
          24184 => x"80", -- $05e78
          24185 => x"80", -- $05e79
          24186 => x"80", -- $05e7a
          24187 => x"80", -- $05e7b
          24188 => x"80", -- $05e7c
          24189 => x"80", -- $05e7d
          24190 => x"80", -- $05e7e
          24191 => x"80", -- $05e7f
          24192 => x"80", -- $05e80
          24193 => x"80", -- $05e81
          24194 => x"7f", -- $05e82
          24195 => x"7f", -- $05e83
          24196 => x"7f", -- $05e84
          24197 => x"7f", -- $05e85
          24198 => x"7f", -- $05e86
          24199 => x"7f", -- $05e87
          24200 => x"7f", -- $05e88
          24201 => x"7f", -- $05e89
          24202 => x"80", -- $05e8a
          24203 => x"80", -- $05e8b
          24204 => x"7f", -- $05e8c
          24205 => x"7f", -- $05e8d
          24206 => x"7f", -- $05e8e
          24207 => x"7f", -- $05e8f
          24208 => x"7f", -- $05e90
          24209 => x"7f", -- $05e91
          24210 => x"7f", -- $05e92
          24211 => x"7f", -- $05e93
          24212 => x"7f", -- $05e94
          24213 => x"7f", -- $05e95
          24214 => x"7f", -- $05e96
          24215 => x"7f", -- $05e97
          24216 => x"7f", -- $05e98
          24217 => x"7f", -- $05e99
          24218 => x"7f", -- $05e9a
          24219 => x"7f", -- $05e9b
          24220 => x"7f", -- $05e9c
          24221 => x"7f", -- $05e9d
          24222 => x"7f", -- $05e9e
          24223 => x"7f", -- $05e9f
          24224 => x"7f", -- $05ea0
          24225 => x"7f", -- $05ea1
          24226 => x"7f", -- $05ea2
          24227 => x"7f", -- $05ea3
          24228 => x"7f", -- $05ea4
          24229 => x"7f", -- $05ea5
          24230 => x"7f", -- $05ea6
          24231 => x"7f", -- $05ea7
          24232 => x"7f", -- $05ea8
          24233 => x"7f", -- $05ea9
          24234 => x"7f", -- $05eaa
          24235 => x"7f", -- $05eab
          24236 => x"7f", -- $05eac
          24237 => x"7f", -- $05ead
          24238 => x"7f", -- $05eae
          24239 => x"7f", -- $05eaf
          24240 => x"7f", -- $05eb0
          24241 => x"7f", -- $05eb1
          24242 => x"7f", -- $05eb2
          24243 => x"7f", -- $05eb3
          24244 => x"7f", -- $05eb4
          24245 => x"7f", -- $05eb5
          24246 => x"7f", -- $05eb6
          24247 => x"7f", -- $05eb7
          24248 => x"7f", -- $05eb8
          24249 => x"7f", -- $05eb9
          24250 => x"7f", -- $05eba
          24251 => x"7f", -- $05ebb
          24252 => x"7f", -- $05ebc
          24253 => x"7f", -- $05ebd
          24254 => x"7f", -- $05ebe
          24255 => x"7f", -- $05ebf
          24256 => x"7f", -- $05ec0
          24257 => x"7f", -- $05ec1
          24258 => x"7f", -- $05ec2
          24259 => x"7f", -- $05ec3
          24260 => x"7f", -- $05ec4
          24261 => x"7f", -- $05ec5
          24262 => x"7f", -- $05ec6
          24263 => x"7f", -- $05ec7
          24264 => x"7f", -- $05ec8
          24265 => x"7f", -- $05ec9
          24266 => x"7f", -- $05eca
          24267 => x"7f", -- $05ecb
          24268 => x"7f", -- $05ecc
          24269 => x"7f", -- $05ecd
          24270 => x"7f", -- $05ece
          24271 => x"7f", -- $05ecf
          24272 => x"7f", -- $05ed0
          24273 => x"7f", -- $05ed1
          24274 => x"7f", -- $05ed2
          24275 => x"7f", -- $05ed3
          24276 => x"7f", -- $05ed4
          24277 => x"7f", -- $05ed5
          24278 => x"7f", -- $05ed6
          24279 => x"7f", -- $05ed7
          24280 => x"7f", -- $05ed8
          24281 => x"7f", -- $05ed9
          24282 => x"7f", -- $05eda
          24283 => x"7f", -- $05edb
          24284 => x"7f", -- $05edc
          24285 => x"7f", -- $05edd
          24286 => x"7f", -- $05ede
          24287 => x"7f", -- $05edf
          24288 => x"7f", -- $05ee0
          24289 => x"7f", -- $05ee1
          24290 => x"7f", -- $05ee2
          24291 => x"7f", -- $05ee3
          24292 => x"7f", -- $05ee4
          24293 => x"7f", -- $05ee5
          24294 => x"7f", -- $05ee6
          24295 => x"7f", -- $05ee7
          24296 => x"7f", -- $05ee8
          24297 => x"7f", -- $05ee9
          24298 => x"7f", -- $05eea
          24299 => x"7f", -- $05eeb
          24300 => x"7f", -- $05eec
          24301 => x"7f", -- $05eed
          24302 => x"7f", -- $05eee
          24303 => x"7f", -- $05eef
          24304 => x"7f", -- $05ef0
          24305 => x"7f", -- $05ef1
          24306 => x"7f", -- $05ef2
          24307 => x"7f", -- $05ef3
          24308 => x"7f", -- $05ef4
          24309 => x"7f", -- $05ef5
          24310 => x"7f", -- $05ef6
          24311 => x"7f", -- $05ef7
          24312 => x"7f", -- $05ef8
          24313 => x"7f", -- $05ef9
          24314 => x"7f", -- $05efa
          24315 => x"7f", -- $05efb
          24316 => x"7f", -- $05efc
          24317 => x"7f", -- $05efd
          24318 => x"7f", -- $05efe
          24319 => x"7f", -- $05eff
          24320 => x"7f", -- $05f00
          24321 => x"7f", -- $05f01
          24322 => x"7f", -- $05f02
          24323 => x"7f", -- $05f03
          24324 => x"7f", -- $05f04
          24325 => x"7f", -- $05f05
          24326 => x"7f", -- $05f06
          24327 => x"7f", -- $05f07
          24328 => x"7f", -- $05f08
          24329 => x"7f", -- $05f09
          24330 => x"7f", -- $05f0a
          24331 => x"7f", -- $05f0b
          24332 => x"7f", -- $05f0c
          24333 => x"7f", -- $05f0d
          24334 => x"7f", -- $05f0e
          24335 => x"7f", -- $05f0f
          24336 => x"7f", -- $05f10
          24337 => x"7f", -- $05f11
          24338 => x"7f", -- $05f12
          24339 => x"7f", -- $05f13
          24340 => x"7f", -- $05f14
          24341 => x"7f", -- $05f15
          24342 => x"7f", -- $05f16
          24343 => x"7f", -- $05f17
          24344 => x"7f", -- $05f18
          24345 => x"80", -- $05f19
          24346 => x"80", -- $05f1a
          24347 => x"80", -- $05f1b
          24348 => x"80", -- $05f1c
          24349 => x"80", -- $05f1d
          24350 => x"80", -- $05f1e
          24351 => x"80", -- $05f1f
          24352 => x"80", -- $05f20
          24353 => x"80", -- $05f21
          24354 => x"7f", -- $05f22
          24355 => x"7f", -- $05f23
          24356 => x"7f", -- $05f24
          24357 => x"80", -- $05f25
          24358 => x"80", -- $05f26
          24359 => x"80", -- $05f27
          24360 => x"80", -- $05f28
          24361 => x"80", -- $05f29
          24362 => x"80", -- $05f2a
          24363 => x"7f", -- $05f2b
          24364 => x"7f", -- $05f2c
          24365 => x"80", -- $05f2d
          24366 => x"80", -- $05f2e
          24367 => x"80", -- $05f2f
          24368 => x"80", -- $05f30
          24369 => x"7f", -- $05f31
          24370 => x"80", -- $05f32
          24371 => x"80", -- $05f33
          24372 => x"80", -- $05f34
          24373 => x"80", -- $05f35
          24374 => x"80", -- $05f36
          24375 => x"80", -- $05f37
          24376 => x"80", -- $05f38
          24377 => x"80", -- $05f39
          24378 => x"80", -- $05f3a
          24379 => x"80", -- $05f3b
          24380 => x"80", -- $05f3c
          24381 => x"80", -- $05f3d
          24382 => x"80", -- $05f3e
          24383 => x"80", -- $05f3f
          24384 => x"80", -- $05f40
          24385 => x"80", -- $05f41
          24386 => x"80", -- $05f42
          24387 => x"80", -- $05f43
          24388 => x"80", -- $05f44
          24389 => x"80", -- $05f45
          24390 => x"80", -- $05f46
          24391 => x"80", -- $05f47
          24392 => x"80", -- $05f48
          24393 => x"80", -- $05f49
          24394 => x"80", -- $05f4a
          24395 => x"80", -- $05f4b
          24396 => x"80", -- $05f4c
          24397 => x"80", -- $05f4d
          24398 => x"80", -- $05f4e
          24399 => x"80", -- $05f4f
          24400 => x"80", -- $05f50
          24401 => x"80", -- $05f51
          24402 => x"80", -- $05f52
          24403 => x"80", -- $05f53
          24404 => x"80", -- $05f54
          24405 => x"80", -- $05f55
          24406 => x"80", -- $05f56
          24407 => x"80", -- $05f57
          24408 => x"80", -- $05f58
          24409 => x"80", -- $05f59
          24410 => x"80", -- $05f5a
          24411 => x"80", -- $05f5b
          24412 => x"80", -- $05f5c
          24413 => x"80", -- $05f5d
          24414 => x"80", -- $05f5e
          24415 => x"80", -- $05f5f
          24416 => x"80", -- $05f60
          24417 => x"80", -- $05f61
          24418 => x"80", -- $05f62
          24419 => x"80", -- $05f63
          24420 => x"80", -- $05f64
          24421 => x"80", -- $05f65
          24422 => x"80", -- $05f66
          24423 => x"80", -- $05f67
          24424 => x"80", -- $05f68
          24425 => x"80", -- $05f69
          24426 => x"80", -- $05f6a
          24427 => x"80", -- $05f6b
          24428 => x"80", -- $05f6c
          24429 => x"80", -- $05f6d
          24430 => x"80", -- $05f6e
          24431 => x"80", -- $05f6f
          24432 => x"80", -- $05f70
          24433 => x"80", -- $05f71
          24434 => x"80", -- $05f72
          24435 => x"80", -- $05f73
          24436 => x"80", -- $05f74
          24437 => x"80", -- $05f75
          24438 => x"80", -- $05f76
          24439 => x"80", -- $05f77
          24440 => x"80", -- $05f78
          24441 => x"80", -- $05f79
          24442 => x"80", -- $05f7a
          24443 => x"80", -- $05f7b
          24444 => x"80", -- $05f7c
          24445 => x"80", -- $05f7d
          24446 => x"80", -- $05f7e
          24447 => x"80", -- $05f7f
          24448 => x"80", -- $05f80
          24449 => x"80", -- $05f81
          24450 => x"80", -- $05f82
          24451 => x"80", -- $05f83
          24452 => x"80", -- $05f84
          24453 => x"80", -- $05f85
          24454 => x"80", -- $05f86
          24455 => x"80", -- $05f87
          24456 => x"80", -- $05f88
          24457 => x"80", -- $05f89
          24458 => x"80", -- $05f8a
          24459 => x"80", -- $05f8b
          24460 => x"80", -- $05f8c
          24461 => x"80", -- $05f8d
          24462 => x"80", -- $05f8e
          24463 => x"80", -- $05f8f
          24464 => x"80", -- $05f90
          24465 => x"80", -- $05f91
          24466 => x"80", -- $05f92
          24467 => x"80", -- $05f93
          24468 => x"80", -- $05f94
          24469 => x"80", -- $05f95
          24470 => x"80", -- $05f96
          24471 => x"80", -- $05f97
          24472 => x"80", -- $05f98
          24473 => x"80", -- $05f99
          24474 => x"80", -- $05f9a
          24475 => x"80", -- $05f9b
          24476 => x"80", -- $05f9c
          24477 => x"80", -- $05f9d
          24478 => x"80", -- $05f9e
          24479 => x"80", -- $05f9f
          24480 => x"80", -- $05fa0
          24481 => x"80", -- $05fa1
          24482 => x"80", -- $05fa2
          24483 => x"80", -- $05fa3
          24484 => x"80", -- $05fa4
          24485 => x"80", -- $05fa5
          24486 => x"80", -- $05fa6
          24487 => x"80", -- $05fa7
          24488 => x"80", -- $05fa8
          24489 => x"80", -- $05fa9
          24490 => x"80", -- $05faa
          24491 => x"80", -- $05fab
          24492 => x"80", -- $05fac
          24493 => x"80", -- $05fad
          24494 => x"80", -- $05fae
          24495 => x"80", -- $05faf
          24496 => x"80", -- $05fb0
          24497 => x"80", -- $05fb1
          24498 => x"80", -- $05fb2
          24499 => x"80", -- $05fb3
          24500 => x"81", -- $05fb4
          24501 => x"80", -- $05fb5
          24502 => x"80", -- $05fb6
          24503 => x"80", -- $05fb7
          24504 => x"81", -- $05fb8
          24505 => x"81", -- $05fb9
          24506 => x"80", -- $05fba
          24507 => x"80", -- $05fbb
          24508 => x"80", -- $05fbc
          24509 => x"80", -- $05fbd
          24510 => x"80", -- $05fbe
          24511 => x"80", -- $05fbf
          24512 => x"80", -- $05fc0
          24513 => x"81", -- $05fc1
          24514 => x"81", -- $05fc2
          24515 => x"81", -- $05fc3
          24516 => x"81", -- $05fc4
          24517 => x"81", -- $05fc5
          24518 => x"81", -- $05fc6
          24519 => x"81", -- $05fc7
          24520 => x"81", -- $05fc8
          24521 => x"81", -- $05fc9
          24522 => x"81", -- $05fca
          24523 => x"81", -- $05fcb
          24524 => x"81", -- $05fcc
          24525 => x"80", -- $05fcd
          24526 => x"81", -- $05fce
          24527 => x"81", -- $05fcf
          24528 => x"81", -- $05fd0
          24529 => x"81", -- $05fd1
          24530 => x"81", -- $05fd2
          24531 => x"81", -- $05fd3
          24532 => x"81", -- $05fd4
          24533 => x"81", -- $05fd5
          24534 => x"81", -- $05fd6
          24535 => x"80", -- $05fd7
          24536 => x"81", -- $05fd8
          24537 => x"81", -- $05fd9
          24538 => x"81", -- $05fda
          24539 => x"80", -- $05fdb
          24540 => x"81", -- $05fdc
          24541 => x"81", -- $05fdd
          24542 => x"81", -- $05fde
          24543 => x"81", -- $05fdf
          24544 => x"81", -- $05fe0
          24545 => x"81", -- $05fe1
          24546 => x"81", -- $05fe2
          24547 => x"80", -- $05fe3
          24548 => x"81", -- $05fe4
          24549 => x"80", -- $05fe5
          24550 => x"80", -- $05fe6
          24551 => x"81", -- $05fe7
          24552 => x"81", -- $05fe8
          24553 => x"81", -- $05fe9
          24554 => x"81", -- $05fea
          24555 => x"81", -- $05feb
          24556 => x"81", -- $05fec
          24557 => x"81", -- $05fed
          24558 => x"81", -- $05fee
          24559 => x"81", -- $05fef
          24560 => x"81", -- $05ff0
          24561 => x"80", -- $05ff1
          24562 => x"80", -- $05ff2
          24563 => x"80", -- $05ff3
          24564 => x"80", -- $05ff4
          24565 => x"80", -- $05ff5
          24566 => x"81", -- $05ff6
          24567 => x"81", -- $05ff7
          24568 => x"80", -- $05ff8
          24569 => x"80", -- $05ff9
          24570 => x"81", -- $05ffa
          24571 => x"81", -- $05ffb
          24572 => x"80", -- $05ffc
          24573 => x"80", -- $05ffd
          24574 => x"80", -- $05ffe
          24575 => x"80", -- $05fff
          24576 => x"80", -- $06000
          24577 => x"80", -- $06001
          24578 => x"81", -- $06002
          24579 => x"81", -- $06003
          24580 => x"81", -- $06004
          24581 => x"81", -- $06005
          24582 => x"81", -- $06006
          24583 => x"81", -- $06007
          24584 => x"81", -- $06008
          24585 => x"81", -- $06009
          24586 => x"81", -- $0600a
          24587 => x"81", -- $0600b
          24588 => x"80", -- $0600c
          24589 => x"81", -- $0600d
          24590 => x"81", -- $0600e
          24591 => x"81", -- $0600f
          24592 => x"81", -- $06010
          24593 => x"81", -- $06011
          24594 => x"80", -- $06012
          24595 => x"81", -- $06013
          24596 => x"80", -- $06014
          24597 => x"80", -- $06015
          24598 => x"81", -- $06016
          24599 => x"80", -- $06017
          24600 => x"80", -- $06018
          24601 => x"80", -- $06019
          24602 => x"80", -- $0601a
          24603 => x"80", -- $0601b
          24604 => x"81", -- $0601c
          24605 => x"80", -- $0601d
          24606 => x"80", -- $0601e
          24607 => x"80", -- $0601f
          24608 => x"80", -- $06020
          24609 => x"81", -- $06021
          24610 => x"81", -- $06022
          24611 => x"81", -- $06023
          24612 => x"81", -- $06024
          24613 => x"81", -- $06025
          24614 => x"80", -- $06026
          24615 => x"81", -- $06027
          24616 => x"81", -- $06028
          24617 => x"81", -- $06029
          24618 => x"81", -- $0602a
          24619 => x"81", -- $0602b
          24620 => x"81", -- $0602c
          24621 => x"81", -- $0602d
          24622 => x"81", -- $0602e
          24623 => x"81", -- $0602f
          24624 => x"81", -- $06030
          24625 => x"81", -- $06031
          24626 => x"81", -- $06032
          24627 => x"80", -- $06033
          24628 => x"80", -- $06034
          24629 => x"80", -- $06035
          24630 => x"80", -- $06036
          24631 => x"80", -- $06037
          24632 => x"80", -- $06038
          24633 => x"81", -- $06039
          24634 => x"81", -- $0603a
          24635 => x"81", -- $0603b
          24636 => x"81", -- $0603c
          24637 => x"80", -- $0603d
          24638 => x"80", -- $0603e
          24639 => x"80", -- $0603f
          24640 => x"80", -- $06040
          24641 => x"80", -- $06041
          24642 => x"80", -- $06042
          24643 => x"80", -- $06043
          24644 => x"80", -- $06044
          24645 => x"80", -- $06045
          24646 => x"80", -- $06046
          24647 => x"80", -- $06047
          24648 => x"80", -- $06048
          24649 => x"80", -- $06049
          24650 => x"80", -- $0604a
          24651 => x"80", -- $0604b
          24652 => x"80", -- $0604c
          24653 => x"80", -- $0604d
          24654 => x"80", -- $0604e
          24655 => x"80", -- $0604f
          24656 => x"80", -- $06050
          24657 => x"80", -- $06051
          24658 => x"80", -- $06052
          24659 => x"80", -- $06053
          24660 => x"80", -- $06054
          24661 => x"80", -- $06055
          24662 => x"80", -- $06056
          24663 => x"80", -- $06057
          24664 => x"80", -- $06058
          24665 => x"80", -- $06059
          24666 => x"80", -- $0605a
          24667 => x"80", -- $0605b
          24668 => x"80", -- $0605c
          24669 => x"80", -- $0605d
          24670 => x"80", -- $0605e
          24671 => x"80", -- $0605f
          24672 => x"80", -- $06060
          24673 => x"80", -- $06061
          24674 => x"80", -- $06062
          24675 => x"80", -- $06063
          24676 => x"80", -- $06064
          24677 => x"80", -- $06065
          24678 => x"80", -- $06066
          24679 => x"80", -- $06067
          24680 => x"80", -- $06068
          24681 => x"80", -- $06069
          24682 => x"80", -- $0606a
          24683 => x"80", -- $0606b
          24684 => x"80", -- $0606c
          24685 => x"80", -- $0606d
          24686 => x"80", -- $0606e
          24687 => x"80", -- $0606f
          24688 => x"80", -- $06070
          24689 => x"80", -- $06071
          24690 => x"80", -- $06072
          24691 => x"80", -- $06073
          24692 => x"80", -- $06074
          24693 => x"80", -- $06075
          24694 => x"80", -- $06076
          24695 => x"80", -- $06077
          24696 => x"80", -- $06078
          24697 => x"80", -- $06079
          24698 => x"81", -- $0607a
          24699 => x"81", -- $0607b
          24700 => x"81", -- $0607c
          24701 => x"81", -- $0607d
          24702 => x"81", -- $0607e
          24703 => x"80", -- $0607f
          24704 => x"80", -- $06080
          24705 => x"80", -- $06081
          24706 => x"80", -- $06082
          24707 => x"80", -- $06083
          24708 => x"80", -- $06084
          24709 => x"81", -- $06085
          24710 => x"81", -- $06086
          24711 => x"81", -- $06087
          24712 => x"81", -- $06088
          24713 => x"81", -- $06089
          24714 => x"81", -- $0608a
          24715 => x"81", -- $0608b
          24716 => x"81", -- $0608c
          24717 => x"81", -- $0608d
          24718 => x"81", -- $0608e
          24719 => x"80", -- $0608f
          24720 => x"81", -- $06090
          24721 => x"80", -- $06091
          24722 => x"81", -- $06092
          24723 => x"81", -- $06093
          24724 => x"81", -- $06094
          24725 => x"81", -- $06095
          24726 => x"81", -- $06096
          24727 => x"81", -- $06097
          24728 => x"81", -- $06098
          24729 => x"81", -- $06099
          24730 => x"81", -- $0609a
          24731 => x"81", -- $0609b
          24732 => x"81", -- $0609c
          24733 => x"81", -- $0609d
          24734 => x"81", -- $0609e
          24735 => x"81", -- $0609f
          24736 => x"81", -- $060a0
          24737 => x"81", -- $060a1
          24738 => x"81", -- $060a2
          24739 => x"81", -- $060a3
          24740 => x"81", -- $060a4
          24741 => x"81", -- $060a5
          24742 => x"81", -- $060a6
          24743 => x"81", -- $060a7
          24744 => x"81", -- $060a8
          24745 => x"81", -- $060a9
          24746 => x"81", -- $060aa
          24747 => x"81", -- $060ab
          24748 => x"81", -- $060ac
          24749 => x"81", -- $060ad
          24750 => x"81", -- $060ae
          24751 => x"81", -- $060af
          24752 => x"81", -- $060b0
          24753 => x"81", -- $060b1
          24754 => x"81", -- $060b2
          24755 => x"81", -- $060b3
          24756 => x"81", -- $060b4
          24757 => x"81", -- $060b5
          24758 => x"81", -- $060b6
          24759 => x"81", -- $060b7
          24760 => x"81", -- $060b8
          24761 => x"81", -- $060b9
          24762 => x"81", -- $060ba
          24763 => x"81", -- $060bb
          24764 => x"81", -- $060bc
          24765 => x"81", -- $060bd
          24766 => x"81", -- $060be
          24767 => x"81", -- $060bf
          24768 => x"81", -- $060c0
          24769 => x"81", -- $060c1
          24770 => x"81", -- $060c2
          24771 => x"81", -- $060c3
          24772 => x"81", -- $060c4
          24773 => x"81", -- $060c5
          24774 => x"81", -- $060c6
          24775 => x"81", -- $060c7
          24776 => x"81", -- $060c8
          24777 => x"81", -- $060c9
          24778 => x"81", -- $060ca
          24779 => x"81", -- $060cb
          24780 => x"81", -- $060cc
          24781 => x"81", -- $060cd
          24782 => x"80", -- $060ce
          24783 => x"80", -- $060cf
          24784 => x"80", -- $060d0
          24785 => x"80", -- $060d1
          24786 => x"80", -- $060d2
          24787 => x"80", -- $060d3
          24788 => x"80", -- $060d4
          24789 => x"80", -- $060d5
          24790 => x"81", -- $060d6
          24791 => x"80", -- $060d7
          24792 => x"80", -- $060d8
          24793 => x"80", -- $060d9
          24794 => x"80", -- $060da
          24795 => x"80", -- $060db
          24796 => x"80", -- $060dc
          24797 => x"80", -- $060dd
          24798 => x"80", -- $060de
          24799 => x"80", -- $060df
          24800 => x"80", -- $060e0
          24801 => x"80", -- $060e1
          24802 => x"80", -- $060e2
          24803 => x"80", -- $060e3
          24804 => x"80", -- $060e4
          24805 => x"80", -- $060e5
          24806 => x"80", -- $060e6
          24807 => x"80", -- $060e7
          24808 => x"80", -- $060e8
          24809 => x"80", -- $060e9
          24810 => x"80", -- $060ea
          24811 => x"80", -- $060eb
          24812 => x"80", -- $060ec
          24813 => x"80", -- $060ed
          24814 => x"80", -- $060ee
          24815 => x"80", -- $060ef
          24816 => x"80", -- $060f0
          24817 => x"80", -- $060f1
          24818 => x"80", -- $060f2
          24819 => x"80", -- $060f3
          24820 => x"80", -- $060f4
          24821 => x"80", -- $060f5
          24822 => x"80", -- $060f6
          24823 => x"80", -- $060f7
          24824 => x"80", -- $060f8
          24825 => x"80", -- $060f9
          24826 => x"80", -- $060fa
          24827 => x"80", -- $060fb
          24828 => x"80", -- $060fc
          24829 => x"80", -- $060fd
          24830 => x"80", -- $060fe
          24831 => x"80", -- $060ff
          24832 => x"80", -- $06100
          24833 => x"80", -- $06101
          24834 => x"80", -- $06102
          24835 => x"80", -- $06103
          24836 => x"80", -- $06104
          24837 => x"80", -- $06105
          24838 => x"80", -- $06106
          24839 => x"80", -- $06107
          24840 => x"80", -- $06108
          24841 => x"80", -- $06109
          24842 => x"80", -- $0610a
          24843 => x"80", -- $0610b
          24844 => x"80", -- $0610c
          24845 => x"80", -- $0610d
          24846 => x"80", -- $0610e
          24847 => x"80", -- $0610f
          24848 => x"80", -- $06110
          24849 => x"80", -- $06111
          24850 => x"80", -- $06112
          24851 => x"80", -- $06113
          24852 => x"80", -- $06114
          24853 => x"80", -- $06115
          24854 => x"80", -- $06116
          24855 => x"80", -- $06117
          24856 => x"80", -- $06118
          24857 => x"80", -- $06119
          24858 => x"7f", -- $0611a
          24859 => x"80", -- $0611b
          24860 => x"80", -- $0611c
          24861 => x"7f", -- $0611d
          24862 => x"7f", -- $0611e
          24863 => x"80", -- $0611f
          24864 => x"80", -- $06120
          24865 => x"80", -- $06121
          24866 => x"7f", -- $06122
          24867 => x"7f", -- $06123
          24868 => x"7f", -- $06124
          24869 => x"7f", -- $06125
          24870 => x"80", -- $06126
          24871 => x"80", -- $06127
          24872 => x"80", -- $06128
          24873 => x"80", -- $06129
          24874 => x"80", -- $0612a
          24875 => x"7f", -- $0612b
          24876 => x"7f", -- $0612c
          24877 => x"7f", -- $0612d
          24878 => x"7f", -- $0612e
          24879 => x"7f", -- $0612f
          24880 => x"7f", -- $06130
          24881 => x"80", -- $06131
          24882 => x"80", -- $06132
          24883 => x"7f", -- $06133
          24884 => x"7f", -- $06134
          24885 => x"7f", -- $06135
          24886 => x"7f", -- $06136
          24887 => x"7f", -- $06137
          24888 => x"7f", -- $06138
          24889 => x"7f", -- $06139
          24890 => x"7f", -- $0613a
          24891 => x"7f", -- $0613b
          24892 => x"7f", -- $0613c
          24893 => x"7f", -- $0613d
          24894 => x"7f", -- $0613e
          24895 => x"7f", -- $0613f
          24896 => x"7f", -- $06140
          24897 => x"7f", -- $06141
          24898 => x"7f", -- $06142
          24899 => x"7f", -- $06143
          24900 => x"7f", -- $06144
          24901 => x"7f", -- $06145
          24902 => x"7f", -- $06146
          24903 => x"7f", -- $06147
          24904 => x"7f", -- $06148
          24905 => x"7f", -- $06149
          24906 => x"7f", -- $0614a
          24907 => x"7f", -- $0614b
          24908 => x"7f", -- $0614c
          24909 => x"7f", -- $0614d
          24910 => x"80", -- $0614e
          24911 => x"7f", -- $0614f
          24912 => x"7f", -- $06150
          24913 => x"80", -- $06151
          24914 => x"7f", -- $06152
          24915 => x"7f", -- $06153
          24916 => x"7f", -- $06154
          24917 => x"7f", -- $06155
          24918 => x"7f", -- $06156
          24919 => x"7f", -- $06157
          24920 => x"80", -- $06158
          24921 => x"80", -- $06159
          24922 => x"80", -- $0615a
          24923 => x"80", -- $0615b
          24924 => x"80", -- $0615c
          24925 => x"80", -- $0615d
          24926 => x"7f", -- $0615e
          24927 => x"80", -- $0615f
          24928 => x"80", -- $06160
          24929 => x"7f", -- $06161
          24930 => x"80", -- $06162
          24931 => x"80", -- $06163
          24932 => x"80", -- $06164
          24933 => x"80", -- $06165
          24934 => x"80", -- $06166
          24935 => x"80", -- $06167
          24936 => x"80", -- $06168
          24937 => x"80", -- $06169
          24938 => x"80", -- $0616a
          24939 => x"80", -- $0616b
          24940 => x"80", -- $0616c
          24941 => x"80", -- $0616d
          24942 => x"80", -- $0616e
          24943 => x"80", -- $0616f
          24944 => x"80", -- $06170
          24945 => x"80", -- $06171
          24946 => x"80", -- $06172
          24947 => x"80", -- $06173
          24948 => x"80", -- $06174
          24949 => x"80", -- $06175
          24950 => x"80", -- $06176
          24951 => x"80", -- $06177
          24952 => x"80", -- $06178
          24953 => x"80", -- $06179
          24954 => x"80", -- $0617a
          24955 => x"80", -- $0617b
          24956 => x"80", -- $0617c
          24957 => x"80", -- $0617d
          24958 => x"80", -- $0617e
          24959 => x"80", -- $0617f
          24960 => x"80", -- $06180
          24961 => x"80", -- $06181
          24962 => x"80", -- $06182
          24963 => x"80", -- $06183
          24964 => x"80", -- $06184
          24965 => x"80", -- $06185
          24966 => x"80", -- $06186
          24967 => x"80", -- $06187
          24968 => x"80", -- $06188
          24969 => x"80", -- $06189
          24970 => x"80", -- $0618a
          24971 => x"80", -- $0618b
          24972 => x"80", -- $0618c
          24973 => x"80", -- $0618d
          24974 => x"80", -- $0618e
          24975 => x"80", -- $0618f
          24976 => x"80", -- $06190
          24977 => x"80", -- $06191
          24978 => x"80", -- $06192
          24979 => x"80", -- $06193
          24980 => x"80", -- $06194
          24981 => x"80", -- $06195
          24982 => x"80", -- $06196
          24983 => x"80", -- $06197
          24984 => x"80", -- $06198
          24985 => x"80", -- $06199
          24986 => x"80", -- $0619a
          24987 => x"80", -- $0619b
          24988 => x"80", -- $0619c
          24989 => x"80", -- $0619d
          24990 => x"80", -- $0619e
          24991 => x"80", -- $0619f
          24992 => x"7f", -- $061a0
          24993 => x"7f", -- $061a1
          24994 => x"7f", -- $061a2
          24995 => x"7f", -- $061a3
          24996 => x"80", -- $061a4
          24997 => x"80", -- $061a5
          24998 => x"80", -- $061a6
          24999 => x"80", -- $061a7
          25000 => x"80", -- $061a8
          25001 => x"7f", -- $061a9
          25002 => x"7f", -- $061aa
          25003 => x"7f", -- $061ab
          25004 => x"7f", -- $061ac
          25005 => x"7f", -- $061ad
          25006 => x"7f", -- $061ae
          25007 => x"7f", -- $061af
          25008 => x"7f", -- $061b0
          25009 => x"7f", -- $061b1
          25010 => x"7f", -- $061b2
          25011 => x"7f", -- $061b3
          25012 => x"7f", -- $061b4
          25013 => x"7f", -- $061b5
          25014 => x"7f", -- $061b6
          25015 => x"7f", -- $061b7
          25016 => x"7f", -- $061b8
          25017 => x"7f", -- $061b9
          25018 => x"7f", -- $061ba
          25019 => x"7f", -- $061bb
          25020 => x"7f", -- $061bc
          25021 => x"7f", -- $061bd
          25022 => x"7f", -- $061be
          25023 => x"7f", -- $061bf
          25024 => x"7f", -- $061c0
          25025 => x"7f", -- $061c1
          25026 => x"7f", -- $061c2
          25027 => x"7f", -- $061c3
          25028 => x"7f", -- $061c4
          25029 => x"7f", -- $061c5
          25030 => x"7f", -- $061c6
          25031 => x"7f", -- $061c7
          25032 => x"7f", -- $061c8
          25033 => x"7f", -- $061c9
          25034 => x"7f", -- $061ca
          25035 => x"7f", -- $061cb
          25036 => x"7f", -- $061cc
          25037 => x"7f", -- $061cd
          25038 => x"7f", -- $061ce
          25039 => x"7f", -- $061cf
          25040 => x"7f", -- $061d0
          25041 => x"7f", -- $061d1
          25042 => x"7f", -- $061d2
          25043 => x"7f", -- $061d3
          25044 => x"7f", -- $061d4
          25045 => x"7f", -- $061d5
          25046 => x"7f", -- $061d6
          25047 => x"7f", -- $061d7
          25048 => x"7f", -- $061d8
          25049 => x"7f", -- $061d9
          25050 => x"7f", -- $061da
          25051 => x"7f", -- $061db
          25052 => x"7f", -- $061dc
          25053 => x"7f", -- $061dd
          25054 => x"7f", -- $061de
          25055 => x"7f", -- $061df
          25056 => x"7f", -- $061e0
          25057 => x"7f", -- $061e1
          25058 => x"7f", -- $061e2
          25059 => x"7f", -- $061e3
          25060 => x"7f", -- $061e4
          25061 => x"7f", -- $061e5
          25062 => x"7f", -- $061e6
          25063 => x"7f", -- $061e7
          25064 => x"7f", -- $061e8
          25065 => x"7f", -- $061e9
          25066 => x"7f", -- $061ea
          25067 => x"7f", -- $061eb
          25068 => x"7f", -- $061ec
          25069 => x"7f", -- $061ed
          25070 => x"7f", -- $061ee
          25071 => x"7f", -- $061ef
          25072 => x"7f", -- $061f0
          25073 => x"7f", -- $061f1
          25074 => x"7f", -- $061f2
          25075 => x"7f", -- $061f3
          25076 => x"7f", -- $061f4
          25077 => x"7f", -- $061f5
          25078 => x"7f", -- $061f6
          25079 => x"7f", -- $061f7
          25080 => x"7f", -- $061f8
          25081 => x"7f", -- $061f9
          25082 => x"7f", -- $061fa
          25083 => x"7f", -- $061fb
          25084 => x"7f", -- $061fc
          25085 => x"7f", -- $061fd
          25086 => x"7f", -- $061fe
          25087 => x"7f", -- $061ff
          25088 => x"7f", -- $06200
          25089 => x"7f", -- $06201
          25090 => x"7f", -- $06202
          25091 => x"7f", -- $06203
          25092 => x"7f", -- $06204
          25093 => x"7f", -- $06205
          25094 => x"7f", -- $06206
          25095 => x"7f", -- $06207
          25096 => x"7f", -- $06208
          25097 => x"7f", -- $06209
          25098 => x"7f", -- $0620a
          25099 => x"7f", -- $0620b
          25100 => x"7f", -- $0620c
          25101 => x"7f", -- $0620d
          25102 => x"7f", -- $0620e
          25103 => x"7f", -- $0620f
          25104 => x"7f", -- $06210
          25105 => x"7f", -- $06211
          25106 => x"7f", -- $06212
          25107 => x"7f", -- $06213
          25108 => x"80", -- $06214
          25109 => x"7f", -- $06215
          25110 => x"7f", -- $06216
          25111 => x"80", -- $06217
          25112 => x"80", -- $06218
          25113 => x"7f", -- $06219
          25114 => x"80", -- $0621a
          25115 => x"80", -- $0621b
          25116 => x"80", -- $0621c
          25117 => x"80", -- $0621d
          25118 => x"80", -- $0621e
          25119 => x"80", -- $0621f
          25120 => x"80", -- $06220
          25121 => x"80", -- $06221
          25122 => x"80", -- $06222
          25123 => x"80", -- $06223
          25124 => x"80", -- $06224
          25125 => x"80", -- $06225
          25126 => x"80", -- $06226
          25127 => x"80", -- $06227
          25128 => x"80", -- $06228
          25129 => x"80", -- $06229
          25130 => x"80", -- $0622a
          25131 => x"80", -- $0622b
          25132 => x"80", -- $0622c
          25133 => x"80", -- $0622d
          25134 => x"80", -- $0622e
          25135 => x"80", -- $0622f
          25136 => x"80", -- $06230
          25137 => x"80", -- $06231
          25138 => x"80", -- $06232
          25139 => x"80", -- $06233
          25140 => x"80", -- $06234
          25141 => x"80", -- $06235
          25142 => x"80", -- $06236
          25143 => x"80", -- $06237
          25144 => x"80", -- $06238
          25145 => x"80", -- $06239
          25146 => x"80", -- $0623a
          25147 => x"80", -- $0623b
          25148 => x"80", -- $0623c
          25149 => x"80", -- $0623d
          25150 => x"80", -- $0623e
          25151 => x"80", -- $0623f
          25152 => x"80", -- $06240
          25153 => x"80", -- $06241
          25154 => x"80", -- $06242
          25155 => x"80", -- $06243
          25156 => x"80", -- $06244
          25157 => x"80", -- $06245
          25158 => x"80", -- $06246
          25159 => x"80", -- $06247
          25160 => x"80", -- $06248
          25161 => x"80", -- $06249
          25162 => x"80", -- $0624a
          25163 => x"80", -- $0624b
          25164 => x"80", -- $0624c
          25165 => x"80", -- $0624d
          25166 => x"80", -- $0624e
          25167 => x"80", -- $0624f
          25168 => x"80", -- $06250
          25169 => x"80", -- $06251
          25170 => x"80", -- $06252
          25171 => x"80", -- $06253
          25172 => x"80", -- $06254
          25173 => x"80", -- $06255
          25174 => x"80", -- $06256
          25175 => x"80", -- $06257
          25176 => x"80", -- $06258
          25177 => x"80", -- $06259
          25178 => x"80", -- $0625a
          25179 => x"80", -- $0625b
          25180 => x"80", -- $0625c
          25181 => x"80", -- $0625d
          25182 => x"80", -- $0625e
          25183 => x"80", -- $0625f
          25184 => x"80", -- $06260
          25185 => x"80", -- $06261
          25186 => x"80", -- $06262
          25187 => x"80", -- $06263
          25188 => x"80", -- $06264
          25189 => x"80", -- $06265
          25190 => x"80", -- $06266
          25191 => x"80", -- $06267
          25192 => x"80", -- $06268
          25193 => x"80", -- $06269
          25194 => x"80", -- $0626a
          25195 => x"80", -- $0626b
          25196 => x"80", -- $0626c
          25197 => x"80", -- $0626d
          25198 => x"80", -- $0626e
          25199 => x"80", -- $0626f
          25200 => x"80", -- $06270
          25201 => x"80", -- $06271
          25202 => x"80", -- $06272
          25203 => x"80", -- $06273
          25204 => x"80", -- $06274
          25205 => x"80", -- $06275
          25206 => x"80", -- $06276
          25207 => x"81", -- $06277
          25208 => x"80", -- $06278
          25209 => x"80", -- $06279
          25210 => x"80", -- $0627a
          25211 => x"81", -- $0627b
          25212 => x"81", -- $0627c
          25213 => x"80", -- $0627d
          25214 => x"80", -- $0627e
          25215 => x"80", -- $0627f
          25216 => x"80", -- $06280
          25217 => x"80", -- $06281
          25218 => x"81", -- $06282
          25219 => x"81", -- $06283
          25220 => x"81", -- $06284
          25221 => x"81", -- $06285
          25222 => x"81", -- $06286
          25223 => x"81", -- $06287
          25224 => x"81", -- $06288
          25225 => x"81", -- $06289
          25226 => x"81", -- $0628a
          25227 => x"81", -- $0628b
          25228 => x"80", -- $0628c
          25229 => x"81", -- $0628d
          25230 => x"81", -- $0628e
          25231 => x"80", -- $0628f
          25232 => x"81", -- $06290
          25233 => x"81", -- $06291
          25234 => x"81", -- $06292
          25235 => x"81", -- $06293
          25236 => x"81", -- $06294
          25237 => x"81", -- $06295
          25238 => x"81", -- $06296
          25239 => x"81", -- $06297
          25240 => x"81", -- $06298
          25241 => x"81", -- $06299
          25242 => x"81", -- $0629a
          25243 => x"81", -- $0629b
          25244 => x"81", -- $0629c
          25245 => x"81", -- $0629d
          25246 => x"81", -- $0629e
          25247 => x"81", -- $0629f
          25248 => x"81", -- $062a0
          25249 => x"81", -- $062a1
          25250 => x"81", -- $062a2
          25251 => x"81", -- $062a3
          25252 => x"81", -- $062a4
          25253 => x"81", -- $062a5
          25254 => x"81", -- $062a6
          25255 => x"81", -- $062a7
          25256 => x"81", -- $062a8
          25257 => x"81", -- $062a9
          25258 => x"81", -- $062aa
          25259 => x"81", -- $062ab
          25260 => x"81", -- $062ac
          25261 => x"81", -- $062ad
          25262 => x"81", -- $062ae
          25263 => x"81", -- $062af
          25264 => x"81", -- $062b0
          25265 => x"81", -- $062b1
          25266 => x"81", -- $062b2
          25267 => x"81", -- $062b3
          25268 => x"81", -- $062b4
          25269 => x"81", -- $062b5
          25270 => x"81", -- $062b6
          25271 => x"81", -- $062b7
          25272 => x"81", -- $062b8
          25273 => x"81", -- $062b9
          25274 => x"81", -- $062ba
          25275 => x"81", -- $062bb
          25276 => x"81", -- $062bc
          25277 => x"81", -- $062bd
          25278 => x"80", -- $062be
          25279 => x"80", -- $062bf
          25280 => x"80", -- $062c0
          25281 => x"80", -- $062c1
          25282 => x"80", -- $062c2
          25283 => x"80", -- $062c3
          25284 => x"80", -- $062c4
          25285 => x"81", -- $062c5
          25286 => x"81", -- $062c6
          25287 => x"81", -- $062c7
          25288 => x"81", -- $062c8
          25289 => x"81", -- $062c9
          25290 => x"80", -- $062ca
          25291 => x"80", -- $062cb
          25292 => x"80", -- $062cc
          25293 => x"80", -- $062cd
          25294 => x"80", -- $062ce
          25295 => x"80", -- $062cf
          25296 => x"80", -- $062d0
          25297 => x"80", -- $062d1
          25298 => x"81", -- $062d2
          25299 => x"81", -- $062d3
          25300 => x"80", -- $062d4
          25301 => x"81", -- $062d5
          25302 => x"81", -- $062d6
          25303 => x"81", -- $062d7
          25304 => x"80", -- $062d8
          25305 => x"80", -- $062d9
          25306 => x"81", -- $062da
          25307 => x"80", -- $062db
          25308 => x"81", -- $062dc
          25309 => x"81", -- $062dd
          25310 => x"81", -- $062de
          25311 => x"81", -- $062df
          25312 => x"81", -- $062e0
          25313 => x"81", -- $062e1
          25314 => x"81", -- $062e2
          25315 => x"81", -- $062e3
          25316 => x"81", -- $062e4
          25317 => x"81", -- $062e5
          25318 => x"80", -- $062e6
          25319 => x"81", -- $062e7
          25320 => x"80", -- $062e8
          25321 => x"81", -- $062e9
          25322 => x"81", -- $062ea
          25323 => x"81", -- $062eb
          25324 => x"81", -- $062ec
          25325 => x"81", -- $062ed
          25326 => x"81", -- $062ee
          25327 => x"81", -- $062ef
          25328 => x"81", -- $062f0
          25329 => x"81", -- $062f1
          25330 => x"81", -- $062f2
          25331 => x"80", -- $062f3
          25332 => x"81", -- $062f4
          25333 => x"81", -- $062f5
          25334 => x"81", -- $062f6
          25335 => x"81", -- $062f7
          25336 => x"81", -- $062f8
          25337 => x"81", -- $062f9
          25338 => x"81", -- $062fa
          25339 => x"81", -- $062fb
          25340 => x"81", -- $062fc
          25341 => x"81", -- $062fd
          25342 => x"81", -- $062fe
          25343 => x"81", -- $062ff
          25344 => x"81", -- $06300
          25345 => x"81", -- $06301
          25346 => x"81", -- $06302
          25347 => x"81", -- $06303
          25348 => x"81", -- $06304
          25349 => x"81", -- $06305
          25350 => x"81", -- $06306
          25351 => x"81", -- $06307
          25352 => x"81", -- $06308
          25353 => x"81", -- $06309
          25354 => x"81", -- $0630a
          25355 => x"81", -- $0630b
          25356 => x"81", -- $0630c
          25357 => x"81", -- $0630d
          25358 => x"81", -- $0630e
          25359 => x"81", -- $0630f
          25360 => x"81", -- $06310
          25361 => x"81", -- $06311
          25362 => x"81", -- $06312
          25363 => x"81", -- $06313
          25364 => x"81", -- $06314
          25365 => x"81", -- $06315
          25366 => x"81", -- $06316
          25367 => x"81", -- $06317
          25368 => x"81", -- $06318
          25369 => x"81", -- $06319
          25370 => x"81", -- $0631a
          25371 => x"81", -- $0631b
          25372 => x"81", -- $0631c
          25373 => x"81", -- $0631d
          25374 => x"81", -- $0631e
          25375 => x"81", -- $0631f
          25376 => x"81", -- $06320
          25377 => x"81", -- $06321
          25378 => x"81", -- $06322
          25379 => x"81", -- $06323
          25380 => x"81", -- $06324
          25381 => x"81", -- $06325
          25382 => x"81", -- $06326
          25383 => x"81", -- $06327
          25384 => x"81", -- $06328
          25385 => x"81", -- $06329
          25386 => x"81", -- $0632a
          25387 => x"81", -- $0632b
          25388 => x"81", -- $0632c
          25389 => x"81", -- $0632d
          25390 => x"81", -- $0632e
          25391 => x"81", -- $0632f
          25392 => x"81", -- $06330
          25393 => x"81", -- $06331
          25394 => x"81", -- $06332
          25395 => x"81", -- $06333
          25396 => x"81", -- $06334
          25397 => x"81", -- $06335
          25398 => x"81", -- $06336
          25399 => x"81", -- $06337
          25400 => x"81", -- $06338
          25401 => x"81", -- $06339
          25402 => x"81", -- $0633a
          25403 => x"81", -- $0633b
          25404 => x"81", -- $0633c
          25405 => x"81", -- $0633d
          25406 => x"81", -- $0633e
          25407 => x"81", -- $0633f
          25408 => x"81", -- $06340
          25409 => x"81", -- $06341
          25410 => x"81", -- $06342
          25411 => x"81", -- $06343
          25412 => x"81", -- $06344
          25413 => x"81", -- $06345
          25414 => x"82", -- $06346
          25415 => x"82", -- $06347
          25416 => x"82", -- $06348
          25417 => x"81", -- $06349
          25418 => x"82", -- $0634a
          25419 => x"82", -- $0634b
          25420 => x"82", -- $0634c
          25421 => x"81", -- $0634d
          25422 => x"81", -- $0634e
          25423 => x"81", -- $0634f
          25424 => x"81", -- $06350
          25425 => x"81", -- $06351
          25426 => x"81", -- $06352
          25427 => x"81", -- $06353
          25428 => x"81", -- $06354
          25429 => x"81", -- $06355
          25430 => x"81", -- $06356
          25431 => x"81", -- $06357
          25432 => x"81", -- $06358
          25433 => x"81", -- $06359
          25434 => x"81", -- $0635a
          25435 => x"81", -- $0635b
          25436 => x"81", -- $0635c
          25437 => x"81", -- $0635d
          25438 => x"81", -- $0635e
          25439 => x"81", -- $0635f
          25440 => x"81", -- $06360
          25441 => x"81", -- $06361
          25442 => x"81", -- $06362
          25443 => x"81", -- $06363
          25444 => x"81", -- $06364
          25445 => x"81", -- $06365
          25446 => x"81", -- $06366
          25447 => x"81", -- $06367
          25448 => x"81", -- $06368
          25449 => x"81", -- $06369
          25450 => x"81", -- $0636a
          25451 => x"81", -- $0636b
          25452 => x"81", -- $0636c
          25453 => x"81", -- $0636d
          25454 => x"81", -- $0636e
          25455 => x"81", -- $0636f
          25456 => x"81", -- $06370
          25457 => x"81", -- $06371
          25458 => x"81", -- $06372
          25459 => x"81", -- $06373
          25460 => x"80", -- $06374
          25461 => x"80", -- $06375
          25462 => x"80", -- $06376
          25463 => x"80", -- $06377
          25464 => x"80", -- $06378
          25465 => x"80", -- $06379
          25466 => x"80", -- $0637a
          25467 => x"80", -- $0637b
          25468 => x"80", -- $0637c
          25469 => x"80", -- $0637d
          25470 => x"80", -- $0637e
          25471 => x"80", -- $0637f
          25472 => x"80", -- $06380
          25473 => x"80", -- $06381
          25474 => x"80", -- $06382
          25475 => x"80", -- $06383
          25476 => x"80", -- $06384
          25477 => x"80", -- $06385
          25478 => x"80", -- $06386
          25479 => x"80", -- $06387
          25480 => x"80", -- $06388
          25481 => x"80", -- $06389
          25482 => x"80", -- $0638a
          25483 => x"80", -- $0638b
          25484 => x"80", -- $0638c
          25485 => x"80", -- $0638d
          25486 => x"80", -- $0638e
          25487 => x"80", -- $0638f
          25488 => x"80", -- $06390
          25489 => x"80", -- $06391
          25490 => x"80", -- $06392
          25491 => x"80", -- $06393
          25492 => x"80", -- $06394
          25493 => x"80", -- $06395
          25494 => x"80", -- $06396
          25495 => x"80", -- $06397
          25496 => x"80", -- $06398
          25497 => x"80", -- $06399
          25498 => x"80", -- $0639a
          25499 => x"80", -- $0639b
          25500 => x"80", -- $0639c
          25501 => x"80", -- $0639d
          25502 => x"80", -- $0639e
          25503 => x"80", -- $0639f
          25504 => x"80", -- $063a0
          25505 => x"80", -- $063a1
          25506 => x"80", -- $063a2
          25507 => x"80", -- $063a3
          25508 => x"80", -- $063a4
          25509 => x"80", -- $063a5
          25510 => x"80", -- $063a6
          25511 => x"80", -- $063a7
          25512 => x"80", -- $063a8
          25513 => x"80", -- $063a9
          25514 => x"80", -- $063aa
          25515 => x"80", -- $063ab
          25516 => x"80", -- $063ac
          25517 => x"80", -- $063ad
          25518 => x"80", -- $063ae
          25519 => x"80", -- $063af
          25520 => x"80", -- $063b0
          25521 => x"80", -- $063b1
          25522 => x"80", -- $063b2
          25523 => x"80", -- $063b3
          25524 => x"80", -- $063b4
          25525 => x"80", -- $063b5
          25526 => x"80", -- $063b6
          25527 => x"80", -- $063b7
          25528 => x"80", -- $063b8
          25529 => x"80", -- $063b9
          25530 => x"80", -- $063ba
          25531 => x"80", -- $063bb
          25532 => x"80", -- $063bc
          25533 => x"80", -- $063bd
          25534 => x"80", -- $063be
          25535 => x"80", -- $063bf
          25536 => x"80", -- $063c0
          25537 => x"80", -- $063c1
          25538 => x"80", -- $063c2
          25539 => x"80", -- $063c3
          25540 => x"80", -- $063c4
          25541 => x"80", -- $063c5
          25542 => x"80", -- $063c6
          25543 => x"80", -- $063c7
          25544 => x"80", -- $063c8
          25545 => x"80", -- $063c9
          25546 => x"80", -- $063ca
          25547 => x"80", -- $063cb
          25548 => x"80", -- $063cc
          25549 => x"80", -- $063cd
          25550 => x"80", -- $063ce
          25551 => x"80", -- $063cf
          25552 => x"80", -- $063d0
          25553 => x"80", -- $063d1
          25554 => x"80", -- $063d2
          25555 => x"80", -- $063d3
          25556 => x"80", -- $063d4
          25557 => x"80", -- $063d5
          25558 => x"80", -- $063d6
          25559 => x"80", -- $063d7
          25560 => x"80", -- $063d8
          25561 => x"80", -- $063d9
          25562 => x"80", -- $063da
          25563 => x"80", -- $063db
          25564 => x"80", -- $063dc
          25565 => x"80", -- $063dd
          25566 => x"80", -- $063de
          25567 => x"80", -- $063df
          25568 => x"80", -- $063e0
          25569 => x"80", -- $063e1
          25570 => x"80", -- $063e2
          25571 => x"80", -- $063e3
          25572 => x"80", -- $063e4
          25573 => x"80", -- $063e5
          25574 => x"80", -- $063e6
          25575 => x"80", -- $063e7
          25576 => x"80", -- $063e8
          25577 => x"80", -- $063e9
          25578 => x"80", -- $063ea
          25579 => x"80", -- $063eb
          25580 => x"80", -- $063ec
          25581 => x"80", -- $063ed
          25582 => x"80", -- $063ee
          25583 => x"80", -- $063ef
          25584 => x"80", -- $063f0
          25585 => x"80", -- $063f1
          25586 => x"80", -- $063f2
          25587 => x"80", -- $063f3
          25588 => x"80", -- $063f4
          25589 => x"80", -- $063f5
          25590 => x"80", -- $063f6
          25591 => x"80", -- $063f7
          25592 => x"80", -- $063f8
          25593 => x"80", -- $063f9
          25594 => x"80", -- $063fa
          25595 => x"80", -- $063fb
          25596 => x"80", -- $063fc
          25597 => x"80", -- $063fd
          25598 => x"80", -- $063fe
          25599 => x"80", -- $063ff
          25600 => x"80", -- $06400
          25601 => x"80", -- $06401
          25602 => x"80", -- $06402
          25603 => x"80", -- $06403
          25604 => x"80", -- $06404
          25605 => x"80", -- $06405
          25606 => x"80", -- $06406
          25607 => x"80", -- $06407
          25608 => x"80", -- $06408
          25609 => x"80", -- $06409
          25610 => x"80", -- $0640a
          25611 => x"80", -- $0640b
          25612 => x"80", -- $0640c
          25613 => x"80", -- $0640d
          25614 => x"80", -- $0640e
          25615 => x"80", -- $0640f
          25616 => x"80", -- $06410
          25617 => x"80", -- $06411
          25618 => x"80", -- $06412
          25619 => x"80", -- $06413
          25620 => x"80", -- $06414
          25621 => x"80", -- $06415
          25622 => x"80", -- $06416
          25623 => x"80", -- $06417
          25624 => x"80", -- $06418
          25625 => x"80", -- $06419
          25626 => x"80", -- $0641a
          25627 => x"80", -- $0641b
          25628 => x"80", -- $0641c
          25629 => x"80", -- $0641d
          25630 => x"80", -- $0641e
          25631 => x"80", -- $0641f
          25632 => x"80", -- $06420
          25633 => x"80", -- $06421
          25634 => x"80", -- $06422
          25635 => x"80", -- $06423
          25636 => x"80", -- $06424
          25637 => x"80", -- $06425
          25638 => x"80", -- $06426
          25639 => x"80", -- $06427
          25640 => x"80", -- $06428
          25641 => x"80", -- $06429
          25642 => x"80", -- $0642a
          25643 => x"80", -- $0642b
          25644 => x"80", -- $0642c
          25645 => x"80", -- $0642d
          25646 => x"80", -- $0642e
          25647 => x"80", -- $0642f
          25648 => x"80", -- $06430
          25649 => x"80", -- $06431
          25650 => x"80", -- $06432
          25651 => x"80", -- $06433
          25652 => x"80", -- $06434
          25653 => x"80", -- $06435
          25654 => x"80", -- $06436
          25655 => x"80", -- $06437
          25656 => x"80", -- $06438
          25657 => x"80", -- $06439
          25658 => x"80", -- $0643a
          25659 => x"80", -- $0643b
          25660 => x"80", -- $0643c
          25661 => x"80", -- $0643d
          25662 => x"80", -- $0643e
          25663 => x"80", -- $0643f
          25664 => x"80", -- $06440
          25665 => x"80", -- $06441
          25666 => x"80", -- $06442
          25667 => x"80", -- $06443
          25668 => x"80", -- $06444
          25669 => x"80", -- $06445
          25670 => x"80", -- $06446
          25671 => x"80", -- $06447
          25672 => x"80", -- $06448
          25673 => x"7f", -- $06449
          25674 => x"7f", -- $0644a
          25675 => x"7f", -- $0644b
          25676 => x"7f", -- $0644c
          25677 => x"7f", -- $0644d
          25678 => x"7f", -- $0644e
          25679 => x"7f", -- $0644f
          25680 => x"7f", -- $06450
          25681 => x"7f", -- $06451
          25682 => x"7f", -- $06452
          25683 => x"7f", -- $06453
          25684 => x"7f", -- $06454
          25685 => x"80", -- $06455
          25686 => x"7f", -- $06456
          25687 => x"7f", -- $06457
          25688 => x"7f", -- $06458
          25689 => x"7f", -- $06459
          25690 => x"7f", -- $0645a
          25691 => x"7f", -- $0645b
          25692 => x"7f", -- $0645c
          25693 => x"7f", -- $0645d
          25694 => x"7f", -- $0645e
          25695 => x"7f", -- $0645f
          25696 => x"7f", -- $06460
          25697 => x"7f", -- $06461
          25698 => x"7f", -- $06462
          25699 => x"7f", -- $06463
          25700 => x"7e", -- $06464
          25701 => x"7e", -- $06465
          25702 => x"7f", -- $06466
          25703 => x"7f", -- $06467
          25704 => x"7f", -- $06468
          25705 => x"7f", -- $06469
          25706 => x"7f", -- $0646a
          25707 => x"7f", -- $0646b
          25708 => x"7f", -- $0646c
          25709 => x"7f", -- $0646d
          25710 => x"7f", -- $0646e
          25711 => x"7f", -- $0646f
          25712 => x"7f", -- $06470
          25713 => x"7f", -- $06471
          25714 => x"7f", -- $06472
          25715 => x"7f", -- $06473
          25716 => x"7f", -- $06474
          25717 => x"7f", -- $06475
          25718 => x"7f", -- $06476
          25719 => x"7f", -- $06477
          25720 => x"7e", -- $06478
          25721 => x"7e", -- $06479
          25722 => x"7e", -- $0647a
          25723 => x"7e", -- $0647b
          25724 => x"7e", -- $0647c
          25725 => x"7e", -- $0647d
          25726 => x"7e", -- $0647e
          25727 => x"7e", -- $0647f
          25728 => x"7f", -- $06480
          25729 => x"7f", -- $06481
          25730 => x"7f", -- $06482
          25731 => x"80", -- $06483
          25732 => x"80", -- $06484
          25733 => x"80", -- $06485
          25734 => x"80", -- $06486
          25735 => x"80", -- $06487
          25736 => x"80", -- $06488
          25737 => x"7f", -- $06489
          25738 => x"7f", -- $0648a
          25739 => x"7f", -- $0648b
          25740 => x"7e", -- $0648c
          25741 => x"7e", -- $0648d
          25742 => x"7e", -- $0648e
          25743 => x"7e", -- $0648f
          25744 => x"7e", -- $06490
          25745 => x"7e", -- $06491
          25746 => x"7e", -- $06492
          25747 => x"7e", -- $06493
          25748 => x"7e", -- $06494
          25749 => x"7f", -- $06495
          25750 => x"7f", -- $06496
          25751 => x"7f", -- $06497
          25752 => x"7f", -- $06498
          25753 => x"80", -- $06499
          25754 => x"80", -- $0649a
          25755 => x"80", -- $0649b
          25756 => x"80", -- $0649c
          25757 => x"7f", -- $0649d
          25758 => x"7f", -- $0649e
          25759 => x"7f", -- $0649f
          25760 => x"7e", -- $064a0
          25761 => x"7e", -- $064a1
          25762 => x"7e", -- $064a2
          25763 => x"7d", -- $064a3
          25764 => x"7d", -- $064a4
          25765 => x"7e", -- $064a5
          25766 => x"7e", -- $064a6
          25767 => x"7e", -- $064a7
          25768 => x"7e", -- $064a8
          25769 => x"7f", -- $064a9
          25770 => x"7f", -- $064aa
          25771 => x"7f", -- $064ab
          25772 => x"7f", -- $064ac
          25773 => x"7f", -- $064ad
          25774 => x"7f", -- $064ae
          25775 => x"7f", -- $064af
          25776 => x"7f", -- $064b0
          25777 => x"7f", -- $064b1
          25778 => x"7e", -- $064b2
          25779 => x"7e", -- $064b3
          25780 => x"7e", -- $064b4
          25781 => x"7e", -- $064b5
          25782 => x"7e", -- $064b6
          25783 => x"7e", -- $064b7
          25784 => x"7e", -- $064b8
          25785 => x"7e", -- $064b9
          25786 => x"7f", -- $064ba
          25787 => x"7f", -- $064bb
          25788 => x"7f", -- $064bc
          25789 => x"7f", -- $064bd
          25790 => x"7f", -- $064be
          25791 => x"7f", -- $064bf
          25792 => x"7f", -- $064c0
          25793 => x"7f", -- $064c1
          25794 => x"7e", -- $064c2
          25795 => x"7e", -- $064c3
          25796 => x"7e", -- $064c4
          25797 => x"7e", -- $064c5
          25798 => x"7e", -- $064c6
          25799 => x"7e", -- $064c7
          25800 => x"7d", -- $064c8
          25801 => x"7d", -- $064c9
          25802 => x"7d", -- $064ca
          25803 => x"7e", -- $064cb
          25804 => x"7e", -- $064cc
          25805 => x"7e", -- $064cd
          25806 => x"7e", -- $064ce
          25807 => x"7f", -- $064cf
          25808 => x"7f", -- $064d0
          25809 => x"7f", -- $064d1
          25810 => x"7f", -- $064d2
          25811 => x"7f", -- $064d3
          25812 => x"7f", -- $064d4
          25813 => x"7f", -- $064d5
          25814 => x"7f", -- $064d6
          25815 => x"7f", -- $064d7
          25816 => x"7f", -- $064d8
          25817 => x"7f", -- $064d9
          25818 => x"7f", -- $064da
          25819 => x"7f", -- $064db
          25820 => x"7f", -- $064dc
          25821 => x"7f", -- $064dd
          25822 => x"7f", -- $064de
          25823 => x"7f", -- $064df
          25824 => x"7f", -- $064e0
          25825 => x"7f", -- $064e1
          25826 => x"7f", -- $064e2
          25827 => x"7f", -- $064e3
          25828 => x"7f", -- $064e4
          25829 => x"7f", -- $064e5
          25830 => x"7f", -- $064e6
          25831 => x"7f", -- $064e7
          25832 => x"7f", -- $064e8
          25833 => x"7f", -- $064e9
          25834 => x"7f", -- $064ea
          25835 => x"7f", -- $064eb
          25836 => x"80", -- $064ec
          25837 => x"80", -- $064ed
          25838 => x"80", -- $064ee
          25839 => x"80", -- $064ef
          25840 => x"80", -- $064f0
          25841 => x"7f", -- $064f1
          25842 => x"7f", -- $064f2
          25843 => x"7f", -- $064f3
          25844 => x"7f", -- $064f4
          25845 => x"7f", -- $064f5
          25846 => x"7f", -- $064f6
          25847 => x"7f", -- $064f7
          25848 => x"7f", -- $064f8
          25849 => x"7f", -- $064f9
          25850 => x"7f", -- $064fa
          25851 => x"7f", -- $064fb
          25852 => x"7f", -- $064fc
          25853 => x"7f", -- $064fd
          25854 => x"7f", -- $064fe
          25855 => x"7f", -- $064ff
          25856 => x"7f", -- $06500
          25857 => x"80", -- $06501
          25858 => x"80", -- $06502
          25859 => x"80", -- $06503
          25860 => x"80", -- $06504
          25861 => x"80", -- $06505
          25862 => x"80", -- $06506
          25863 => x"80", -- $06507
          25864 => x"80", -- $06508
          25865 => x"80", -- $06509
          25866 => x"80", -- $0650a
          25867 => x"80", -- $0650b
          25868 => x"80", -- $0650c
          25869 => x"80", -- $0650d
          25870 => x"80", -- $0650e
          25871 => x"80", -- $0650f
          25872 => x"80", -- $06510
          25873 => x"80", -- $06511
          25874 => x"80", -- $06512
          25875 => x"80", -- $06513
          25876 => x"80", -- $06514
          25877 => x"80", -- $06515
          25878 => x"80", -- $06516
          25879 => x"80", -- $06517
          25880 => x"80", -- $06518
          25881 => x"80", -- $06519
          25882 => x"80", -- $0651a
          25883 => x"80", -- $0651b
          25884 => x"80", -- $0651c
          25885 => x"80", -- $0651d
          25886 => x"80", -- $0651e
          25887 => x"80", -- $0651f
          25888 => x"80", -- $06520
          25889 => x"80", -- $06521
          25890 => x"80", -- $06522
          25891 => x"80", -- $06523
          25892 => x"80", -- $06524
          25893 => x"80", -- $06525
          25894 => x"80", -- $06526
          25895 => x"80", -- $06527
          25896 => x"80", -- $06528
          25897 => x"80", -- $06529
          25898 => x"80", -- $0652a
          25899 => x"80", -- $0652b
          25900 => x"80", -- $0652c
          25901 => x"80", -- $0652d
          25902 => x"80", -- $0652e
          25903 => x"80", -- $0652f
          25904 => x"80", -- $06530
          25905 => x"80", -- $06531
          25906 => x"80", -- $06532
          25907 => x"80", -- $06533
          25908 => x"80", -- $06534
          25909 => x"80", -- $06535
          25910 => x"80", -- $06536
          25911 => x"80", -- $06537
          25912 => x"80", -- $06538
          25913 => x"80", -- $06539
          25914 => x"80", -- $0653a
          25915 => x"80", -- $0653b
          25916 => x"80", -- $0653c
          25917 => x"80", -- $0653d
          25918 => x"80", -- $0653e
          25919 => x"80", -- $0653f
          25920 => x"80", -- $06540
          25921 => x"80", -- $06541
          25922 => x"80", -- $06542
          25923 => x"80", -- $06543
          25924 => x"80", -- $06544
          25925 => x"80", -- $06545
          25926 => x"80", -- $06546
          25927 => x"80", -- $06547
          25928 => x"80", -- $06548
          25929 => x"80", -- $06549
          25930 => x"80", -- $0654a
          25931 => x"80", -- $0654b
          25932 => x"80", -- $0654c
          25933 => x"80", -- $0654d
          25934 => x"80", -- $0654e
          25935 => x"80", -- $0654f
          25936 => x"80", -- $06550
          25937 => x"80", -- $06551
          25938 => x"80", -- $06552
          25939 => x"80", -- $06553
          25940 => x"80", -- $06554
          25941 => x"80", -- $06555
          25942 => x"80", -- $06556
          25943 => x"80", -- $06557
          25944 => x"80", -- $06558
          25945 => x"80", -- $06559
          25946 => x"80", -- $0655a
          25947 => x"80", -- $0655b
          25948 => x"80", -- $0655c
          25949 => x"80", -- $0655d
          25950 => x"80", -- $0655e
          25951 => x"80", -- $0655f
          25952 => x"80", -- $06560
          25953 => x"80", -- $06561
          25954 => x"80", -- $06562
          25955 => x"80", -- $06563
          25956 => x"80", -- $06564
          25957 => x"80", -- $06565
          25958 => x"80", -- $06566
          25959 => x"80", -- $06567
          25960 => x"80", -- $06568
          25961 => x"80", -- $06569
          25962 => x"80", -- $0656a
          25963 => x"80", -- $0656b
          25964 => x"80", -- $0656c
          25965 => x"80", -- $0656d
          25966 => x"80", -- $0656e
          25967 => x"80", -- $0656f
          25968 => x"80", -- $06570
          25969 => x"80", -- $06571
          25970 => x"80", -- $06572
          25971 => x"80", -- $06573
          25972 => x"80", -- $06574
          25973 => x"80", -- $06575
          25974 => x"80", -- $06576
          25975 => x"80", -- $06577
          25976 => x"80", -- $06578
          25977 => x"80", -- $06579
          25978 => x"80", -- $0657a
          25979 => x"80", -- $0657b
          25980 => x"80", -- $0657c
          25981 => x"80", -- $0657d
          25982 => x"80", -- $0657e
          25983 => x"80", -- $0657f
          25984 => x"80", -- $06580
          25985 => x"80", -- $06581
          25986 => x"80", -- $06582
          25987 => x"80", -- $06583
          25988 => x"80", -- $06584
          25989 => x"80", -- $06585
          25990 => x"80", -- $06586
          25991 => x"80", -- $06587
          25992 => x"80", -- $06588
          25993 => x"80", -- $06589
          25994 => x"80", -- $0658a
          25995 => x"80", -- $0658b
          25996 => x"80", -- $0658c
          25997 => x"80", -- $0658d
          25998 => x"80", -- $0658e
          25999 => x"80", -- $0658f
          26000 => x"80", -- $06590
          26001 => x"80", -- $06591
          26002 => x"80", -- $06592
          26003 => x"80", -- $06593
          26004 => x"80", -- $06594
          26005 => x"80", -- $06595
          26006 => x"80", -- $06596
          26007 => x"80", -- $06597
          26008 => x"80", -- $06598
          26009 => x"80", -- $06599
          26010 => x"80", -- $0659a
          26011 => x"80", -- $0659b
          26012 => x"80", -- $0659c
          26013 => x"80", -- $0659d
          26014 => x"80", -- $0659e
          26015 => x"80", -- $0659f
          26016 => x"80", -- $065a0
          26017 => x"80", -- $065a1
          26018 => x"80", -- $065a2
          26019 => x"80", -- $065a3
          26020 => x"80", -- $065a4
          26021 => x"80", -- $065a5
          26022 => x"80", -- $065a6
          26023 => x"80", -- $065a7
          26024 => x"80", -- $065a8
          26025 => x"80", -- $065a9
          26026 => x"80", -- $065aa
          26027 => x"80", -- $065ab
          26028 => x"80", -- $065ac
          26029 => x"81", -- $065ad
          26030 => x"80", -- $065ae
          26031 => x"81", -- $065af
          26032 => x"81", -- $065b0
          26033 => x"80", -- $065b1
          26034 => x"80", -- $065b2
          26035 => x"80", -- $065b3
          26036 => x"80", -- $065b4
          26037 => x"80", -- $065b5
          26038 => x"80", -- $065b6
          26039 => x"80", -- $065b7
          26040 => x"80", -- $065b8
          26041 => x"80", -- $065b9
          26042 => x"80", -- $065ba
          26043 => x"80", -- $065bb
          26044 => x"80", -- $065bc
          26045 => x"81", -- $065bd
          26046 => x"81", -- $065be
          26047 => x"81", -- $065bf
          26048 => x"81", -- $065c0
          26049 => x"80", -- $065c1
          26050 => x"80", -- $065c2
          26051 => x"80", -- $065c3
          26052 => x"80", -- $065c4
          26053 => x"80", -- $065c5
          26054 => x"81", -- $065c6
          26055 => x"81", -- $065c7
          26056 => x"81", -- $065c8
          26057 => x"81", -- $065c9
          26058 => x"81", -- $065ca
          26059 => x"81", -- $065cb
          26060 => x"81", -- $065cc
          26061 => x"81", -- $065cd
          26062 => x"80", -- $065ce
          26063 => x"80", -- $065cf
          26064 => x"80", -- $065d0
          26065 => x"80", -- $065d1
          26066 => x"80", -- $065d2
          26067 => x"80", -- $065d3
          26068 => x"80", -- $065d4
          26069 => x"80", -- $065d5
          26070 => x"80", -- $065d6
          26071 => x"80", -- $065d7
          26072 => x"80", -- $065d8
          26073 => x"80", -- $065d9
          26074 => x"80", -- $065da
          26075 => x"80", -- $065db
          26076 => x"80", -- $065dc
          26077 => x"80", -- $065dd
          26078 => x"80", -- $065de
          26079 => x"80", -- $065df
          26080 => x"80", -- $065e0
          26081 => x"80", -- $065e1
          26082 => x"80", -- $065e2
          26083 => x"80", -- $065e3
          26084 => x"80", -- $065e4
          26085 => x"80", -- $065e5
          26086 => x"80", -- $065e6
          26087 => x"80", -- $065e7
          26088 => x"80", -- $065e8
          26089 => x"80", -- $065e9
          26090 => x"80", -- $065ea
          26091 => x"80", -- $065eb
          26092 => x"80", -- $065ec
          26093 => x"80", -- $065ed
          26094 => x"80", -- $065ee
          26095 => x"80", -- $065ef
          26096 => x"80", -- $065f0
          26097 => x"80", -- $065f1
          26098 => x"80", -- $065f2
          26099 => x"80", -- $065f3
          26100 => x"80", -- $065f4
          26101 => x"80", -- $065f5
          26102 => x"80", -- $065f6
          26103 => x"80", -- $065f7
          26104 => x"80", -- $065f8
          26105 => x"80", -- $065f9
          26106 => x"80", -- $065fa
          26107 => x"80", -- $065fb
          26108 => x"80", -- $065fc
          26109 => x"80", -- $065fd
          26110 => x"80", -- $065fe
          26111 => x"80", -- $065ff
          26112 => x"80", -- $06600
          26113 => x"80", -- $06601
          26114 => x"80", -- $06602
          26115 => x"80", -- $06603
          26116 => x"80", -- $06604
          26117 => x"80", -- $06605
          26118 => x"80", -- $06606
          26119 => x"80", -- $06607
          26120 => x"80", -- $06608
          26121 => x"80", -- $06609
          26122 => x"80", -- $0660a
          26123 => x"80", -- $0660b
          26124 => x"80", -- $0660c
          26125 => x"80", -- $0660d
          26126 => x"80", -- $0660e
          26127 => x"80", -- $0660f
          26128 => x"80", -- $06610
          26129 => x"80", -- $06611
          26130 => x"80", -- $06612
          26131 => x"80", -- $06613
          26132 => x"80", -- $06614
          26133 => x"80", -- $06615
          26134 => x"80", -- $06616
          26135 => x"80", -- $06617
          26136 => x"80", -- $06618
          26137 => x"80", -- $06619
          26138 => x"80", -- $0661a
          26139 => x"80", -- $0661b
          26140 => x"80", -- $0661c
          26141 => x"80", -- $0661d
          26142 => x"80", -- $0661e
          26143 => x"80", -- $0661f
          26144 => x"80", -- $06620
          26145 => x"80", -- $06621
          26146 => x"80", -- $06622
          26147 => x"80", -- $06623
          26148 => x"80", -- $06624
          26149 => x"80", -- $06625
          26150 => x"80", -- $06626
          26151 => x"80", -- $06627
          26152 => x"80", -- $06628
          26153 => x"80", -- $06629
          26154 => x"80", -- $0662a
          26155 => x"80", -- $0662b
          26156 => x"80", -- $0662c
          26157 => x"80", -- $0662d
          26158 => x"80", -- $0662e
          26159 => x"80", -- $0662f
          26160 => x"80", -- $06630
          26161 => x"80", -- $06631
          26162 => x"80", -- $06632
          26163 => x"80", -- $06633
          26164 => x"80", -- $06634
          26165 => x"80", -- $06635
          26166 => x"80", -- $06636
          26167 => x"80", -- $06637
          26168 => x"80", -- $06638
          26169 => x"80", -- $06639
          26170 => x"80", -- $0663a
          26171 => x"80", -- $0663b
          26172 => x"81", -- $0663c
          26173 => x"81", -- $0663d
          26174 => x"81", -- $0663e
          26175 => x"81", -- $0663f
          26176 => x"81", -- $06640
          26177 => x"81", -- $06641
          26178 => x"81", -- $06642
          26179 => x"81", -- $06643
          26180 => x"81", -- $06644
          26181 => x"81", -- $06645
          26182 => x"81", -- $06646
          26183 => x"81", -- $06647
          26184 => x"81", -- $06648
          26185 => x"81", -- $06649
          26186 => x"81", -- $0664a
          26187 => x"81", -- $0664b
          26188 => x"82", -- $0664c
          26189 => x"82", -- $0664d
          26190 => x"82", -- $0664e
          26191 => x"81", -- $0664f
          26192 => x"82", -- $06650
          26193 => x"82", -- $06651
          26194 => x"82", -- $06652
          26195 => x"82", -- $06653
          26196 => x"82", -- $06654
          26197 => x"82", -- $06655
          26198 => x"82", -- $06656
          26199 => x"82", -- $06657
          26200 => x"82", -- $06658
          26201 => x"82", -- $06659
          26202 => x"82", -- $0665a
          26203 => x"82", -- $0665b
          26204 => x"82", -- $0665c
          26205 => x"82", -- $0665d
          26206 => x"82", -- $0665e
          26207 => x"82", -- $0665f
          26208 => x"82", -- $06660
          26209 => x"82", -- $06661
          26210 => x"82", -- $06662
          26211 => x"82", -- $06663
          26212 => x"82", -- $06664
          26213 => x"82", -- $06665
          26214 => x"82", -- $06666
          26215 => x"82", -- $06667
          26216 => x"82", -- $06668
          26217 => x"82", -- $06669
          26218 => x"82", -- $0666a
          26219 => x"81", -- $0666b
          26220 => x"82", -- $0666c
          26221 => x"82", -- $0666d
          26222 => x"82", -- $0666e
          26223 => x"81", -- $0666f
          26224 => x"81", -- $06670
          26225 => x"82", -- $06671
          26226 => x"81", -- $06672
          26227 => x"82", -- $06673
          26228 => x"81", -- $06674
          26229 => x"81", -- $06675
          26230 => x"81", -- $06676
          26231 => x"81", -- $06677
          26232 => x"81", -- $06678
          26233 => x"81", -- $06679
          26234 => x"81", -- $0667a
          26235 => x"81", -- $0667b
          26236 => x"81", -- $0667c
          26237 => x"81", -- $0667d
          26238 => x"81", -- $0667e
          26239 => x"81", -- $0667f
          26240 => x"81", -- $06680
          26241 => x"81", -- $06681
          26242 => x"81", -- $06682
          26243 => x"81", -- $06683
          26244 => x"81", -- $06684
          26245 => x"81", -- $06685
          26246 => x"81", -- $06686
          26247 => x"81", -- $06687
          26248 => x"81", -- $06688
          26249 => x"81", -- $06689
          26250 => x"81", -- $0668a
          26251 => x"81", -- $0668b
          26252 => x"81", -- $0668c
          26253 => x"81", -- $0668d
          26254 => x"81", -- $0668e
          26255 => x"81", -- $0668f
          26256 => x"81", -- $06690
          26257 => x"81", -- $06691
          26258 => x"81", -- $06692
          26259 => x"81", -- $06693
          26260 => x"81", -- $06694
          26261 => x"81", -- $06695
          26262 => x"81", -- $06696
          26263 => x"81", -- $06697
          26264 => x"81", -- $06698
          26265 => x"81", -- $06699
          26266 => x"81", -- $0669a
          26267 => x"81", -- $0669b
          26268 => x"81", -- $0669c
          26269 => x"81", -- $0669d
          26270 => x"80", -- $0669e
          26271 => x"80", -- $0669f
          26272 => x"80", -- $066a0
          26273 => x"80", -- $066a1
          26274 => x"80", -- $066a2
          26275 => x"80", -- $066a3
          26276 => x"80", -- $066a4
          26277 => x"80", -- $066a5
          26278 => x"80", -- $066a6
          26279 => x"80", -- $066a7
          26280 => x"80", -- $066a8
          26281 => x"80", -- $066a9
          26282 => x"80", -- $066aa
          26283 => x"80", -- $066ab
          26284 => x"80", -- $066ac
          26285 => x"80", -- $066ad
          26286 => x"80", -- $066ae
          26287 => x"80", -- $066af
          26288 => x"80", -- $066b0
          26289 => x"80", -- $066b1
          26290 => x"80", -- $066b2
          26291 => x"80", -- $066b3
          26292 => x"80", -- $066b4
          26293 => x"80", -- $066b5
          26294 => x"80", -- $066b6
          26295 => x"80", -- $066b7
          26296 => x"80", -- $066b8
          26297 => x"80", -- $066b9
          26298 => x"80", -- $066ba
          26299 => x"80", -- $066bb
          26300 => x"80", -- $066bc
          26301 => x"80", -- $066bd
          26302 => x"80", -- $066be
          26303 => x"80", -- $066bf
          26304 => x"80", -- $066c0
          26305 => x"80", -- $066c1
          26306 => x"80", -- $066c2
          26307 => x"80", -- $066c3
          26308 => x"80", -- $066c4
          26309 => x"80", -- $066c5
          26310 => x"80", -- $066c6
          26311 => x"80", -- $066c7
          26312 => x"80", -- $066c8
          26313 => x"80", -- $066c9
          26314 => x"80", -- $066ca
          26315 => x"80", -- $066cb
          26316 => x"80", -- $066cc
          26317 => x"80", -- $066cd
          26318 => x"80", -- $066ce
          26319 => x"80", -- $066cf
          26320 => x"80", -- $066d0
          26321 => x"80", -- $066d1
          26322 => x"80", -- $066d2
          26323 => x"80", -- $066d3
          26324 => x"80", -- $066d4
          26325 => x"80", -- $066d5
          26326 => x"80", -- $066d6
          26327 => x"80", -- $066d7
          26328 => x"80", -- $066d8
          26329 => x"80", -- $066d9
          26330 => x"80", -- $066da
          26331 => x"80", -- $066db
          26332 => x"80", -- $066dc
          26333 => x"80", -- $066dd
          26334 => x"80", -- $066de
          26335 => x"80", -- $066df
          26336 => x"80", -- $066e0
          26337 => x"80", -- $066e1
          26338 => x"80", -- $066e2
          26339 => x"80", -- $066e3
          26340 => x"80", -- $066e4
          26341 => x"80", -- $066e5
          26342 => x"80", -- $066e6
          26343 => x"80", -- $066e7
          26344 => x"80", -- $066e8
          26345 => x"80", -- $066e9
          26346 => x"80", -- $066ea
          26347 => x"80", -- $066eb
          26348 => x"80", -- $066ec
          26349 => x"80", -- $066ed
          26350 => x"80", -- $066ee
          26351 => x"80", -- $066ef
          26352 => x"80", -- $066f0
          26353 => x"80", -- $066f1
          26354 => x"80", -- $066f2
          26355 => x"80", -- $066f3
          26356 => x"80", -- $066f4
          26357 => x"80", -- $066f5
          26358 => x"80", -- $066f6
          26359 => x"80", -- $066f7
          26360 => x"80", -- $066f8
          26361 => x"80", -- $066f9
          26362 => x"80", -- $066fa
          26363 => x"80", -- $066fb
          26364 => x"80", -- $066fc
          26365 => x"80", -- $066fd
          26366 => x"80", -- $066fe
          26367 => x"80", -- $066ff
          26368 => x"80", -- $06700
          26369 => x"80", -- $06701
          26370 => x"80", -- $06702
          26371 => x"80", -- $06703
          26372 => x"80", -- $06704
          26373 => x"7f", -- $06705
          26374 => x"80", -- $06706
          26375 => x"80", -- $06707
          26376 => x"80", -- $06708
          26377 => x"80", -- $06709
          26378 => x"80", -- $0670a
          26379 => x"80", -- $0670b
          26380 => x"80", -- $0670c
          26381 => x"80", -- $0670d
          26382 => x"80", -- $0670e
          26383 => x"80", -- $0670f
          26384 => x"80", -- $06710
          26385 => x"80", -- $06711
          26386 => x"80", -- $06712
          26387 => x"80", -- $06713
          26388 => x"80", -- $06714
          26389 => x"80", -- $06715
          26390 => x"80", -- $06716
          26391 => x"80", -- $06717
          26392 => x"80", -- $06718
          26393 => x"80", -- $06719
          26394 => x"80", -- $0671a
          26395 => x"80", -- $0671b
          26396 => x"80", -- $0671c
          26397 => x"80", -- $0671d
          26398 => x"80", -- $0671e
          26399 => x"80", -- $0671f
          26400 => x"80", -- $06720
          26401 => x"80", -- $06721
          26402 => x"80", -- $06722
          26403 => x"80", -- $06723
          26404 => x"80", -- $06724
          26405 => x"80", -- $06725
          26406 => x"80", -- $06726
          26407 => x"80", -- $06727
          26408 => x"80", -- $06728
          26409 => x"80", -- $06729
          26410 => x"80", -- $0672a
          26411 => x"80", -- $0672b
          26412 => x"80", -- $0672c
          26413 => x"80", -- $0672d
          26414 => x"80", -- $0672e
          26415 => x"80", -- $0672f
          26416 => x"80", -- $06730
          26417 => x"80", -- $06731
          26418 => x"80", -- $06732
          26419 => x"80", -- $06733
          26420 => x"80", -- $06734
          26421 => x"80", -- $06735
          26422 => x"80", -- $06736
          26423 => x"80", -- $06737
          26424 => x"80", -- $06738
          26425 => x"80", -- $06739
          26426 => x"80", -- $0673a
          26427 => x"80", -- $0673b
          26428 => x"80", -- $0673c
          26429 => x"80", -- $0673d
          26430 => x"80", -- $0673e
          26431 => x"80", -- $0673f
          26432 => x"80", -- $06740
          26433 => x"80", -- $06741
          26434 => x"80", -- $06742
          26435 => x"80", -- $06743
          26436 => x"80", -- $06744
          26437 => x"80", -- $06745
          26438 => x"80", -- $06746
          26439 => x"80", -- $06747
          26440 => x"80", -- $06748
          26441 => x"80", -- $06749
          26442 => x"80", -- $0674a
          26443 => x"80", -- $0674b
          26444 => x"80", -- $0674c
          26445 => x"80", -- $0674d
          26446 => x"80", -- $0674e
          26447 => x"80", -- $0674f
          26448 => x"80", -- $06750
          26449 => x"80", -- $06751
          26450 => x"80", -- $06752
          26451 => x"80", -- $06753
          26452 => x"80", -- $06754
          26453 => x"80", -- $06755
          26454 => x"80", -- $06756
          26455 => x"80", -- $06757
          26456 => x"80", -- $06758
          26457 => x"80", -- $06759
          26458 => x"80", -- $0675a
          26459 => x"80", -- $0675b
          26460 => x"80", -- $0675c
          26461 => x"80", -- $0675d
          26462 => x"80", -- $0675e
          26463 => x"80", -- $0675f
          26464 => x"80", -- $06760
          26465 => x"80", -- $06761
          26466 => x"80", -- $06762
          26467 => x"80", -- $06763
          26468 => x"80", -- $06764
          26469 => x"80", -- $06765
          26470 => x"80", -- $06766
          26471 => x"80", -- $06767
          26472 => x"80", -- $06768
          26473 => x"80", -- $06769
          26474 => x"80", -- $0676a
          26475 => x"80", -- $0676b
          26476 => x"80", -- $0676c
          26477 => x"7f", -- $0676d
          26478 => x"7f", -- $0676e
          26479 => x"7f", -- $0676f
          26480 => x"7f", -- $06770
          26481 => x"7f", -- $06771
          26482 => x"7f", -- $06772
          26483 => x"7f", -- $06773
          26484 => x"7f", -- $06774
          26485 => x"7f", -- $06775
          26486 => x"7f", -- $06776
          26487 => x"7f", -- $06777
          26488 => x"7f", -- $06778
          26489 => x"80", -- $06779
          26490 => x"7f", -- $0677a
          26491 => x"80", -- $0677b
          26492 => x"7f", -- $0677c
          26493 => x"7f", -- $0677d
          26494 => x"7f", -- $0677e
          26495 => x"7f", -- $0677f
          26496 => x"7f", -- $06780
          26497 => x"7f", -- $06781
          26498 => x"7f", -- $06782
          26499 => x"7f", -- $06783
          26500 => x"7f", -- $06784
          26501 => x"7f", -- $06785
          26502 => x"7f", -- $06786
          26503 => x"7f", -- $06787
          26504 => x"7f", -- $06788
          26505 => x"7f", -- $06789
          26506 => x"7f", -- $0678a
          26507 => x"7f", -- $0678b
          26508 => x"7f", -- $0678c
          26509 => x"7f", -- $0678d
          26510 => x"7f", -- $0678e
          26511 => x"7f", -- $0678f
          26512 => x"7f", -- $06790
          26513 => x"7f", -- $06791
          26514 => x"7f", -- $06792
          26515 => x"7f", -- $06793
          26516 => x"7f", -- $06794
          26517 => x"7f", -- $06795
          26518 => x"7f", -- $06796
          26519 => x"7f", -- $06797
          26520 => x"7f", -- $06798
          26521 => x"7f", -- $06799
          26522 => x"7f", -- $0679a
          26523 => x"7f", -- $0679b
          26524 => x"7f", -- $0679c
          26525 => x"7f", -- $0679d
          26526 => x"7f", -- $0679e
          26527 => x"7f", -- $0679f
          26528 => x"7f", -- $067a0
          26529 => x"7f", -- $067a1
          26530 => x"7f", -- $067a2
          26531 => x"7f", -- $067a3
          26532 => x"7f", -- $067a4
          26533 => x"7f", -- $067a5
          26534 => x"7e", -- $067a6
          26535 => x"7e", -- $067a7
          26536 => x"7e", -- $067a8
          26537 => x"7f", -- $067a9
          26538 => x"7f", -- $067aa
          26539 => x"7f", -- $067ab
          26540 => x"7f", -- $067ac
          26541 => x"7e", -- $067ad
          26542 => x"7e", -- $067ae
          26543 => x"7e", -- $067af
          26544 => x"7e", -- $067b0
          26545 => x"7e", -- $067b1
          26546 => x"7e", -- $067b2
          26547 => x"7e", -- $067b3
          26548 => x"7e", -- $067b4
          26549 => x"7e", -- $067b5
          26550 => x"7e", -- $067b6
          26551 => x"7e", -- $067b7
          26552 => x"7e", -- $067b8
          26553 => x"7e", -- $067b9
          26554 => x"7e", -- $067ba
          26555 => x"7e", -- $067bb
          26556 => x"7e", -- $067bc
          26557 => x"7e", -- $067bd
          26558 => x"7e", -- $067be
          26559 => x"7e", -- $067bf
          26560 => x"7e", -- $067c0
          26561 => x"7e", -- $067c1
          26562 => x"7e", -- $067c2
          26563 => x"7e", -- $067c3
          26564 => x"7e", -- $067c4
          26565 => x"7e", -- $067c5
          26566 => x"7e", -- $067c6
          26567 => x"7d", -- $067c7
          26568 => x"7d", -- $067c8
          26569 => x"7d", -- $067c9
          26570 => x"7d", -- $067ca
          26571 => x"7d", -- $067cb
          26572 => x"7d", -- $067cc
          26573 => x"7d", -- $067cd
          26574 => x"7d", -- $067ce
          26575 => x"7d", -- $067cf
          26576 => x"7d", -- $067d0
          26577 => x"7d", -- $067d1
          26578 => x"7d", -- $067d2
          26579 => x"7d", -- $067d3
          26580 => x"7d", -- $067d4
          26581 => x"7d", -- $067d5
          26582 => x"7d", -- $067d6
          26583 => x"7d", -- $067d7
          26584 => x"7d", -- $067d8
          26585 => x"7d", -- $067d9
          26586 => x"7d", -- $067da
          26587 => x"7d", -- $067db
          26588 => x"7d", -- $067dc
          26589 => x"7d", -- $067dd
          26590 => x"7d", -- $067de
          26591 => x"7d", -- $067df
          26592 => x"7d", -- $067e0
          26593 => x"7d", -- $067e1
          26594 => x"7d", -- $067e2
          26595 => x"7d", -- $067e3
          26596 => x"7d", -- $067e4
          26597 => x"7d", -- $067e5
          26598 => x"7d", -- $067e6
          26599 => x"7d", -- $067e7
          26600 => x"7d", -- $067e8
          26601 => x"7d", -- $067e9
          26602 => x"7e", -- $067ea
          26603 => x"7d", -- $067eb
          26604 => x"7e", -- $067ec
          26605 => x"7e", -- $067ed
          26606 => x"7e", -- $067ee
          26607 => x"7e", -- $067ef
          26608 => x"7e", -- $067f0
          26609 => x"7e", -- $067f1
          26610 => x"7e", -- $067f2
          26611 => x"7e", -- $067f3
          26612 => x"7e", -- $067f4
          26613 => x"7e", -- $067f5
          26614 => x"7e", -- $067f6
          26615 => x"7e", -- $067f7
          26616 => x"7e", -- $067f8
          26617 => x"7e", -- $067f9
          26618 => x"7e", -- $067fa
          26619 => x"7e", -- $067fb
          26620 => x"7e", -- $067fc
          26621 => x"7e", -- $067fd
          26622 => x"7e", -- $067fe
          26623 => x"7e", -- $067ff
          26624 => x"7e", -- $06800
          26625 => x"7e", -- $06801
          26626 => x"7e", -- $06802
          26627 => x"7e", -- $06803
          26628 => x"7e", -- $06804
          26629 => x"7e", -- $06805
          26630 => x"7e", -- $06806
          26631 => x"7f", -- $06807
          26632 => x"7f", -- $06808
          26633 => x"7f", -- $06809
          26634 => x"7f", -- $0680a
          26635 => x"7f", -- $0680b
          26636 => x"7f", -- $0680c
          26637 => x"7f", -- $0680d
          26638 => x"7f", -- $0680e
          26639 => x"7f", -- $0680f
          26640 => x"7f", -- $06810
          26641 => x"7f", -- $06811
          26642 => x"7f", -- $06812
          26643 => x"7f", -- $06813
          26644 => x"7f", -- $06814
          26645 => x"7f", -- $06815
          26646 => x"7f", -- $06816
          26647 => x"7f", -- $06817
          26648 => x"7f", -- $06818
          26649 => x"7f", -- $06819
          26650 => x"7f", -- $0681a
          26651 => x"7f", -- $0681b
          26652 => x"7f", -- $0681c
          26653 => x"7f", -- $0681d
          26654 => x"7f", -- $0681e
          26655 => x"7f", -- $0681f
          26656 => x"7f", -- $06820
          26657 => x"7f", -- $06821
          26658 => x"7f", -- $06822
          26659 => x"7f", -- $06823
          26660 => x"7f", -- $06824
          26661 => x"7f", -- $06825
          26662 => x"7f", -- $06826
          26663 => x"7f", -- $06827
          26664 => x"7f", -- $06828
          26665 => x"7f", -- $06829
          26666 => x"7f", -- $0682a
          26667 => x"7f", -- $0682b
          26668 => x"7f", -- $0682c
          26669 => x"7f", -- $0682d
          26670 => x"7f", -- $0682e
          26671 => x"7f", -- $0682f
          26672 => x"80", -- $06830
          26673 => x"80", -- $06831
          26674 => x"7f", -- $06832
          26675 => x"7f", -- $06833
          26676 => x"7f", -- $06834
          26677 => x"7f", -- $06835
          26678 => x"7f", -- $06836
          26679 => x"7f", -- $06837
          26680 => x"80", -- $06838
          26681 => x"80", -- $06839
          26682 => x"80", -- $0683a
          26683 => x"80", -- $0683b
          26684 => x"80", -- $0683c
          26685 => x"80", -- $0683d
          26686 => x"80", -- $0683e
          26687 => x"80", -- $0683f
          26688 => x"80", -- $06840
          26689 => x"80", -- $06841
          26690 => x"80", -- $06842
          26691 => x"80", -- $06843
          26692 => x"80", -- $06844
          26693 => x"80", -- $06845
          26694 => x"80", -- $06846
          26695 => x"80", -- $06847
          26696 => x"80", -- $06848
          26697 => x"80", -- $06849
          26698 => x"80", -- $0684a
          26699 => x"80", -- $0684b
          26700 => x"80", -- $0684c
          26701 => x"80", -- $0684d
          26702 => x"80", -- $0684e
          26703 => x"80", -- $0684f
          26704 => x"80", -- $06850
          26705 => x"80", -- $06851
          26706 => x"80", -- $06852
          26707 => x"80", -- $06853
          26708 => x"80", -- $06854
          26709 => x"80", -- $06855
          26710 => x"80", -- $06856
          26711 => x"80", -- $06857
          26712 => x"80", -- $06858
          26713 => x"80", -- $06859
          26714 => x"80", -- $0685a
          26715 => x"80", -- $0685b
          26716 => x"80", -- $0685c
          26717 => x"80", -- $0685d
          26718 => x"80", -- $0685e
          26719 => x"80", -- $0685f
          26720 => x"80", -- $06860
          26721 => x"80", -- $06861
          26722 => x"80", -- $06862
          26723 => x"80", -- $06863
          26724 => x"80", -- $06864
          26725 => x"80", -- $06865
          26726 => x"80", -- $06866
          26727 => x"80", -- $06867
          26728 => x"80", -- $06868
          26729 => x"80", -- $06869
          26730 => x"80", -- $0686a
          26731 => x"80", -- $0686b
          26732 => x"80", -- $0686c
          26733 => x"80", -- $0686d
          26734 => x"80", -- $0686e
          26735 => x"80", -- $0686f
          26736 => x"80", -- $06870
          26737 => x"80", -- $06871
          26738 => x"80", -- $06872
          26739 => x"80", -- $06873
          26740 => x"80", -- $06874
          26741 => x"80", -- $06875
          26742 => x"80", -- $06876
          26743 => x"80", -- $06877
          26744 => x"80", -- $06878
          26745 => x"80", -- $06879
          26746 => x"80", -- $0687a
          26747 => x"80", -- $0687b
          26748 => x"80", -- $0687c
          26749 => x"80", -- $0687d
          26750 => x"80", -- $0687e
          26751 => x"80", -- $0687f
          26752 => x"80", -- $06880
          26753 => x"80", -- $06881
          26754 => x"80", -- $06882
          26755 => x"80", -- $06883
          26756 => x"80", -- $06884
          26757 => x"80", -- $06885
          26758 => x"80", -- $06886
          26759 => x"80", -- $06887
          26760 => x"80", -- $06888
          26761 => x"80", -- $06889
          26762 => x"80", -- $0688a
          26763 => x"80", -- $0688b
          26764 => x"80", -- $0688c
          26765 => x"80", -- $0688d
          26766 => x"80", -- $0688e
          26767 => x"80", -- $0688f
          26768 => x"80", -- $06890
          26769 => x"80", -- $06891
          26770 => x"80", -- $06892
          26771 => x"80", -- $06893
          26772 => x"80", -- $06894
          26773 => x"80", -- $06895
          26774 => x"80", -- $06896
          26775 => x"80", -- $06897
          26776 => x"80", -- $06898
          26777 => x"80", -- $06899
          26778 => x"80", -- $0689a
          26779 => x"80", -- $0689b
          26780 => x"80", -- $0689c
          26781 => x"80", -- $0689d
          26782 => x"80", -- $0689e
          26783 => x"80", -- $0689f
          26784 => x"80", -- $068a0
          26785 => x"80", -- $068a1
          26786 => x"80", -- $068a2
          26787 => x"80", -- $068a3
          26788 => x"80", -- $068a4
          26789 => x"80", -- $068a5
          26790 => x"80", -- $068a6
          26791 => x"80", -- $068a7
          26792 => x"80", -- $068a8
          26793 => x"80", -- $068a9
          26794 => x"80", -- $068aa
          26795 => x"80", -- $068ab
          26796 => x"80", -- $068ac
          26797 => x"80", -- $068ad
          26798 => x"80", -- $068ae
          26799 => x"80", -- $068af
          26800 => x"80", -- $068b0
          26801 => x"80", -- $068b1
          26802 => x"80", -- $068b2
          26803 => x"80", -- $068b3
          26804 => x"80", -- $068b4
          26805 => x"80", -- $068b5
          26806 => x"80", -- $068b6
          26807 => x"80", -- $068b7
          26808 => x"80", -- $068b8
          26809 => x"80", -- $068b9
          26810 => x"80", -- $068ba
          26811 => x"80", -- $068bb
          26812 => x"80", -- $068bc
          26813 => x"80", -- $068bd
          26814 => x"80", -- $068be
          26815 => x"80", -- $068bf
          26816 => x"80", -- $068c0
          26817 => x"80", -- $068c1
          26818 => x"80", -- $068c2
          26819 => x"80", -- $068c3
          26820 => x"80", -- $068c4
          26821 => x"80", -- $068c5
          26822 => x"81", -- $068c6
          26823 => x"81", -- $068c7
          26824 => x"81", -- $068c8
          26825 => x"81", -- $068c9
          26826 => x"81", -- $068ca
          26827 => x"81", -- $068cb
          26828 => x"81", -- $068cc
          26829 => x"81", -- $068cd
          26830 => x"81", -- $068ce
          26831 => x"81", -- $068cf
          26832 => x"81", -- $068d0
          26833 => x"81", -- $068d1
          26834 => x"81", -- $068d2
          26835 => x"81", -- $068d3
          26836 => x"81", -- $068d4
          26837 => x"81", -- $068d5
          26838 => x"81", -- $068d6
          26839 => x"81", -- $068d7
          26840 => x"81", -- $068d8
          26841 => x"81", -- $068d9
          26842 => x"81", -- $068da
          26843 => x"81", -- $068db
          26844 => x"81", -- $068dc
          26845 => x"82", -- $068dd
          26846 => x"82", -- $068de
          26847 => x"82", -- $068df
          26848 => x"82", -- $068e0
          26849 => x"82", -- $068e1
          26850 => x"82", -- $068e2
          26851 => x"82", -- $068e3
          26852 => x"82", -- $068e4
          26853 => x"82", -- $068e5
          26854 => x"82", -- $068e6
          26855 => x"82", -- $068e7
          26856 => x"82", -- $068e8
          26857 => x"82", -- $068e9
          26858 => x"82", -- $068ea
          26859 => x"82", -- $068eb
          26860 => x"82", -- $068ec
          26861 => x"82", -- $068ed
          26862 => x"82", -- $068ee
          26863 => x"82", -- $068ef
          26864 => x"82", -- $068f0
          26865 => x"82", -- $068f1
          26866 => x"82", -- $068f2
          26867 => x"82", -- $068f3
          26868 => x"82", -- $068f4
          26869 => x"82", -- $068f5
          26870 => x"82", -- $068f6
          26871 => x"82", -- $068f7
          26872 => x"82", -- $068f8
          26873 => x"82", -- $068f9
          26874 => x"82", -- $068fa
          26875 => x"82", -- $068fb
          26876 => x"82", -- $068fc
          26877 => x"82", -- $068fd
          26878 => x"82", -- $068fe
          26879 => x"82", -- $068ff
          26880 => x"82", -- $06900
          26881 => x"82", -- $06901
          26882 => x"82", -- $06902
          26883 => x"82", -- $06903
          26884 => x"82", -- $06904
          26885 => x"82", -- $06905
          26886 => x"82", -- $06906
          26887 => x"82", -- $06907
          26888 => x"82", -- $06908
          26889 => x"83", -- $06909
          26890 => x"83", -- $0690a
          26891 => x"83", -- $0690b
          26892 => x"83", -- $0690c
          26893 => x"83", -- $0690d
          26894 => x"83", -- $0690e
          26895 => x"83", -- $0690f
          26896 => x"83", -- $06910
          26897 => x"83", -- $06911
          26898 => x"83", -- $06912
          26899 => x"83", -- $06913
          26900 => x"83", -- $06914
          26901 => x"83", -- $06915
          26902 => x"83", -- $06916
          26903 => x"83", -- $06917
          26904 => x"83", -- $06918
          26905 => x"83", -- $06919
          26906 => x"83", -- $0691a
          26907 => x"83", -- $0691b
          26908 => x"83", -- $0691c
          26909 => x"83", -- $0691d
          26910 => x"83", -- $0691e
          26911 => x"83", -- $0691f
          26912 => x"83", -- $06920
          26913 => x"83", -- $06921
          26914 => x"83", -- $06922
          26915 => x"83", -- $06923
          26916 => x"83", -- $06924
          26917 => x"83", -- $06925
          26918 => x"83", -- $06926
          26919 => x"83", -- $06927
          26920 => x"83", -- $06928
          26921 => x"83", -- $06929
          26922 => x"83", -- $0692a
          26923 => x"83", -- $0692b
          26924 => x"83", -- $0692c
          26925 => x"83", -- $0692d
          26926 => x"83", -- $0692e
          26927 => x"83", -- $0692f
          26928 => x"83", -- $06930
          26929 => x"83", -- $06931
          26930 => x"83", -- $06932
          26931 => x"83", -- $06933
          26932 => x"84", -- $06934
          26933 => x"83", -- $06935
          26934 => x"84", -- $06936
          26935 => x"83", -- $06937
          26936 => x"83", -- $06938
          26937 => x"83", -- $06939
          26938 => x"84", -- $0693a
          26939 => x"83", -- $0693b
          26940 => x"83", -- $0693c
          26941 => x"83", -- $0693d
          26942 => x"83", -- $0693e
          26943 => x"83", -- $0693f
          26944 => x"83", -- $06940
          26945 => x"83", -- $06941
          26946 => x"83", -- $06942
          26947 => x"83", -- $06943
          26948 => x"83", -- $06944
          26949 => x"83", -- $06945
          26950 => x"83", -- $06946
          26951 => x"83", -- $06947
          26952 => x"83", -- $06948
          26953 => x"83", -- $06949
          26954 => x"83", -- $0694a
          26955 => x"83", -- $0694b
          26956 => x"83", -- $0694c
          26957 => x"83", -- $0694d
          26958 => x"83", -- $0694e
          26959 => x"83", -- $0694f
          26960 => x"83", -- $06950
          26961 => x"83", -- $06951
          26962 => x"83", -- $06952
          26963 => x"83", -- $06953
          26964 => x"83", -- $06954
          26965 => x"83", -- $06955
          26966 => x"83", -- $06956
          26967 => x"83", -- $06957
          26968 => x"83", -- $06958
          26969 => x"83", -- $06959
          26970 => x"83", -- $0695a
          26971 => x"83", -- $0695b
          26972 => x"83", -- $0695c
          26973 => x"83", -- $0695d
          26974 => x"83", -- $0695e
          26975 => x"83", -- $0695f
          26976 => x"83", -- $06960
          26977 => x"83", -- $06961
          26978 => x"83", -- $06962
          26979 => x"83", -- $06963
          26980 => x"83", -- $06964
          26981 => x"83", -- $06965
          26982 => x"83", -- $06966
          26983 => x"83", -- $06967
          26984 => x"83", -- $06968
          26985 => x"83", -- $06969
          26986 => x"83", -- $0696a
          26987 => x"83", -- $0696b
          26988 => x"83", -- $0696c
          26989 => x"83", -- $0696d
          26990 => x"83", -- $0696e
          26991 => x"83", -- $0696f
          26992 => x"83", -- $06970
          26993 => x"83", -- $06971
          26994 => x"83", -- $06972
          26995 => x"83", -- $06973
          26996 => x"83", -- $06974
          26997 => x"83", -- $06975
          26998 => x"83", -- $06976
          26999 => x"83", -- $06977
          27000 => x"83", -- $06978
          27001 => x"83", -- $06979
          27002 => x"83", -- $0697a
          27003 => x"83", -- $0697b
          27004 => x"82", -- $0697c
          27005 => x"82", -- $0697d
          27006 => x"82", -- $0697e
          27007 => x"82", -- $0697f
          27008 => x"82", -- $06980
          27009 => x"82", -- $06981
          27010 => x"82", -- $06982
          27011 => x"82", -- $06983
          27012 => x"82", -- $06984
          27013 => x"82", -- $06985
          27014 => x"82", -- $06986
          27015 => x"82", -- $06987
          27016 => x"82", -- $06988
          27017 => x"82", -- $06989
          27018 => x"82", -- $0698a
          27019 => x"82", -- $0698b
          27020 => x"82", -- $0698c
          27021 => x"82", -- $0698d
          27022 => x"82", -- $0698e
          27023 => x"82", -- $0698f
          27024 => x"82", -- $06990
          27025 => x"82", -- $06991
          27026 => x"82", -- $06992
          27027 => x"82", -- $06993
          27028 => x"82", -- $06994
          27029 => x"82", -- $06995
          27030 => x"82", -- $06996
          27031 => x"82", -- $06997
          27032 => x"82", -- $06998
          27033 => x"82", -- $06999
          27034 => x"82", -- $0699a
          27035 => x"82", -- $0699b
          27036 => x"82", -- $0699c
          27037 => x"82", -- $0699d
          27038 => x"82", -- $0699e
          27039 => x"82", -- $0699f
          27040 => x"82", -- $069a0
          27041 => x"82", -- $069a1
          27042 => x"82", -- $069a2
          27043 => x"82", -- $069a3
          27044 => x"82", -- $069a4
          27045 => x"82", -- $069a5
          27046 => x"82", -- $069a6
          27047 => x"82", -- $069a7
          27048 => x"82", -- $069a8
          27049 => x"82", -- $069a9
          27050 => x"82", -- $069aa
          27051 => x"82", -- $069ab
          27052 => x"82", -- $069ac
          27053 => x"82", -- $069ad
          27054 => x"82", -- $069ae
          27055 => x"82", -- $069af
          27056 => x"81", -- $069b0
          27057 => x"81", -- $069b1
          27058 => x"82", -- $069b2
          27059 => x"81", -- $069b3
          27060 => x"81", -- $069b4
          27061 => x"81", -- $069b5
          27062 => x"81", -- $069b6
          27063 => x"82", -- $069b7
          27064 => x"82", -- $069b8
          27065 => x"81", -- $069b9
          27066 => x"81", -- $069ba
          27067 => x"81", -- $069bb
          27068 => x"81", -- $069bc
          27069 => x"81", -- $069bd
          27070 => x"81", -- $069be
          27071 => x"81", -- $069bf
          27072 => x"81", -- $069c0
          27073 => x"81", -- $069c1
          27074 => x"81", -- $069c2
          27075 => x"81", -- $069c3
          27076 => x"81", -- $069c4
          27077 => x"81", -- $069c5
          27078 => x"81", -- $069c6
          27079 => x"81", -- $069c7
          27080 => x"81", -- $069c8
          27081 => x"81", -- $069c9
          27082 => x"81", -- $069ca
          27083 => x"81", -- $069cb
          27084 => x"81", -- $069cc
          27085 => x"81", -- $069cd
          27086 => x"81", -- $069ce
          27087 => x"81", -- $069cf
          27088 => x"81", -- $069d0
          27089 => x"81", -- $069d1
          27090 => x"81", -- $069d2
          27091 => x"81", -- $069d3
          27092 => x"81", -- $069d4
          27093 => x"81", -- $069d5
          27094 => x"81", -- $069d6
          27095 => x"81", -- $069d7
          27096 => x"81", -- $069d8
          27097 => x"81", -- $069d9
          27098 => x"81", -- $069da
          27099 => x"81", -- $069db
          27100 => x"81", -- $069dc
          27101 => x"81", -- $069dd
          27102 => x"81", -- $069de
          27103 => x"81", -- $069df
          27104 => x"81", -- $069e0
          27105 => x"81", -- $069e1
          27106 => x"81", -- $069e2
          27107 => x"81", -- $069e3
          27108 => x"81", -- $069e4
          27109 => x"81", -- $069e5
          27110 => x"81", -- $069e6
          27111 => x"81", -- $069e7
          27112 => x"81", -- $069e8
          27113 => x"81", -- $069e9
          27114 => x"81", -- $069ea
          27115 => x"81", -- $069eb
          27116 => x"81", -- $069ec
          27117 => x"81", -- $069ed
          27118 => x"81", -- $069ee
          27119 => x"81", -- $069ef
          27120 => x"81", -- $069f0
          27121 => x"81", -- $069f1
          27122 => x"81", -- $069f2
          27123 => x"80", -- $069f3
          27124 => x"81", -- $069f4
          27125 => x"81", -- $069f5
          27126 => x"81", -- $069f6
          27127 => x"81", -- $069f7
          27128 => x"81", -- $069f8
          27129 => x"81", -- $069f9
          27130 => x"81", -- $069fa
          27131 => x"81", -- $069fb
          27132 => x"81", -- $069fc
          27133 => x"80", -- $069fd
          27134 => x"80", -- $069fe
          27135 => x"80", -- $069ff
          27136 => x"80", -- $06a00
          27137 => x"80", -- $06a01
          27138 => x"80", -- $06a02
          27139 => x"80", -- $06a03
          27140 => x"80", -- $06a04
          27141 => x"80", -- $06a05
          27142 => x"80", -- $06a06
          27143 => x"80", -- $06a07
          27144 => x"80", -- $06a08
          27145 => x"80", -- $06a09
          27146 => x"80", -- $06a0a
          27147 => x"80", -- $06a0b
          27148 => x"80", -- $06a0c
          27149 => x"80", -- $06a0d
          27150 => x"80", -- $06a0e
          27151 => x"80", -- $06a0f
          27152 => x"80", -- $06a10
          27153 => x"80", -- $06a11
          27154 => x"80", -- $06a12
          27155 => x"80", -- $06a13
          27156 => x"80", -- $06a14
          27157 => x"80", -- $06a15
          27158 => x"80", -- $06a16
          27159 => x"80", -- $06a17
          27160 => x"80", -- $06a18
          27161 => x"80", -- $06a19
          27162 => x"80", -- $06a1a
          27163 => x"80", -- $06a1b
          27164 => x"80", -- $06a1c
          27165 => x"80", -- $06a1d
          27166 => x"80", -- $06a1e
          27167 => x"80", -- $06a1f
          27168 => x"80", -- $06a20
          27169 => x"80", -- $06a21
          27170 => x"80", -- $06a22
          27171 => x"80", -- $06a23
          27172 => x"80", -- $06a24
          27173 => x"80", -- $06a25
          27174 => x"80", -- $06a26
          27175 => x"80", -- $06a27
          27176 => x"80", -- $06a28
          27177 => x"80", -- $06a29
          27178 => x"80", -- $06a2a
          27179 => x"80", -- $06a2b
          27180 => x"80", -- $06a2c
          27181 => x"80", -- $06a2d
          27182 => x"80", -- $06a2e
          27183 => x"80", -- $06a2f
          27184 => x"80", -- $06a30
          27185 => x"80", -- $06a31
          27186 => x"80", -- $06a32
          27187 => x"80", -- $06a33
          27188 => x"80", -- $06a34
          27189 => x"80", -- $06a35
          27190 => x"80", -- $06a36
          27191 => x"80", -- $06a37
          27192 => x"80", -- $06a38
          27193 => x"7f", -- $06a39
          27194 => x"7f", -- $06a3a
          27195 => x"7f", -- $06a3b
          27196 => x"7f", -- $06a3c
          27197 => x"7f", -- $06a3d
          27198 => x"7f", -- $06a3e
          27199 => x"7f", -- $06a3f
          27200 => x"7f", -- $06a40
          27201 => x"7f", -- $06a41
          27202 => x"7f", -- $06a42
          27203 => x"7f", -- $06a43
          27204 => x"7f", -- $06a44
          27205 => x"7f", -- $06a45
          27206 => x"7f", -- $06a46
          27207 => x"7f", -- $06a47
          27208 => x"7f", -- $06a48
          27209 => x"7f", -- $06a49
          27210 => x"7e", -- $06a4a
          27211 => x"7e", -- $06a4b
          27212 => x"7e", -- $06a4c
          27213 => x"7e", -- $06a4d
          27214 => x"7e", -- $06a4e
          27215 => x"7e", -- $06a4f
          27216 => x"7e", -- $06a50
          27217 => x"7e", -- $06a51
          27218 => x"7e", -- $06a52
          27219 => x"7e", -- $06a53
          27220 => x"7e", -- $06a54
          27221 => x"7e", -- $06a55
          27222 => x"7e", -- $06a56
          27223 => x"7e", -- $06a57
          27224 => x"7e", -- $06a58
          27225 => x"7e", -- $06a59
          27226 => x"7e", -- $06a5a
          27227 => x"7e", -- $06a5b
          27228 => x"7e", -- $06a5c
          27229 => x"7e", -- $06a5d
          27230 => x"7e", -- $06a5e
          27231 => x"7e", -- $06a5f
          27232 => x"7e", -- $06a60
          27233 => x"7e", -- $06a61
          27234 => x"7e", -- $06a62
          27235 => x"7e", -- $06a63
          27236 => x"7e", -- $06a64
          27237 => x"7e", -- $06a65
          27238 => x"7e", -- $06a66
          27239 => x"7e", -- $06a67
          27240 => x"7e", -- $06a68
          27241 => x"7e", -- $06a69
          27242 => x"7e", -- $06a6a
          27243 => x"7e", -- $06a6b
          27244 => x"7e", -- $06a6c
          27245 => x"7e", -- $06a6d
          27246 => x"7e", -- $06a6e
          27247 => x"7e", -- $06a6f
          27248 => x"7e", -- $06a70
          27249 => x"7e", -- $06a71
          27250 => x"7e", -- $06a72
          27251 => x"7e", -- $06a73
          27252 => x"7e", -- $06a74
          27253 => x"7e", -- $06a75
          27254 => x"7e", -- $06a76
          27255 => x"7e", -- $06a77
          27256 => x"7e", -- $06a78
          27257 => x"7e", -- $06a79
          27258 => x"7e", -- $06a7a
          27259 => x"7e", -- $06a7b
          27260 => x"7e", -- $06a7c
          27261 => x"7e", -- $06a7d
          27262 => x"7e", -- $06a7e
          27263 => x"7e", -- $06a7f
          27264 => x"7e", -- $06a80
          27265 => x"7e", -- $06a81
          27266 => x"7e", -- $06a82
          27267 => x"7e", -- $06a83
          27268 => x"7e", -- $06a84
          27269 => x"7e", -- $06a85
          27270 => x"7e", -- $06a86
          27271 => x"7e", -- $06a87
          27272 => x"7e", -- $06a88
          27273 => x"7e", -- $06a89
          27274 => x"7e", -- $06a8a
          27275 => x"7e", -- $06a8b
          27276 => x"7e", -- $06a8c
          27277 => x"7e", -- $06a8d
          27278 => x"7e", -- $06a8e
          27279 => x"7e", -- $06a8f
          27280 => x"7e", -- $06a90
          27281 => x"7e", -- $06a91
          27282 => x"7e", -- $06a92
          27283 => x"7e", -- $06a93
          27284 => x"7e", -- $06a94
          27285 => x"7e", -- $06a95
          27286 => x"7e", -- $06a96
          27287 => x"7e", -- $06a97
          27288 => x"7e", -- $06a98
          27289 => x"7e", -- $06a99
          27290 => x"7e", -- $06a9a
          27291 => x"7e", -- $06a9b
          27292 => x"7e", -- $06a9c
          27293 => x"7e", -- $06a9d
          27294 => x"7e", -- $06a9e
          27295 => x"7e", -- $06a9f
          27296 => x"7e", -- $06aa0
          27297 => x"7e", -- $06aa1
          27298 => x"7e", -- $06aa2
          27299 => x"7e", -- $06aa3
          27300 => x"7e", -- $06aa4
          27301 => x"7e", -- $06aa5
          27302 => x"7e", -- $06aa6
          27303 => x"7d", -- $06aa7
          27304 => x"7d", -- $06aa8
          27305 => x"7d", -- $06aa9
          27306 => x"7d", -- $06aaa
          27307 => x"7e", -- $06aab
          27308 => x"7e", -- $06aac
          27309 => x"7e", -- $06aad
          27310 => x"7e", -- $06aae
          27311 => x"7e", -- $06aaf
          27312 => x"7e", -- $06ab0
          27313 => x"7d", -- $06ab1
          27314 => x"7d", -- $06ab2
          27315 => x"7d", -- $06ab3
          27316 => x"7d", -- $06ab4
          27317 => x"7d", -- $06ab5
          27318 => x"7d", -- $06ab6
          27319 => x"7d", -- $06ab7
          27320 => x"7d", -- $06ab8
          27321 => x"7d", -- $06ab9
          27322 => x"7d", -- $06aba
          27323 => x"7d", -- $06abb
          27324 => x"7d", -- $06abc
          27325 => x"7d", -- $06abd
          27326 => x"7d", -- $06abe
          27327 => x"7d", -- $06abf
          27328 => x"7d", -- $06ac0
          27329 => x"7d", -- $06ac1
          27330 => x"7d", -- $06ac2
          27331 => x"7d", -- $06ac3
          27332 => x"7d", -- $06ac4
          27333 => x"7d", -- $06ac5
          27334 => x"7d", -- $06ac6
          27335 => x"7d", -- $06ac7
          27336 => x"7d", -- $06ac8
          27337 => x"7d", -- $06ac9
          27338 => x"7d", -- $06aca
          27339 => x"7d", -- $06acb
          27340 => x"7d", -- $06acc
          27341 => x"7d", -- $06acd
          27342 => x"7c", -- $06ace
          27343 => x"7c", -- $06acf
          27344 => x"7c", -- $06ad0
          27345 => x"7c", -- $06ad1
          27346 => x"7d", -- $06ad2
          27347 => x"7d", -- $06ad3
          27348 => x"7d", -- $06ad4
          27349 => x"7d", -- $06ad5
          27350 => x"7d", -- $06ad6
          27351 => x"7c", -- $06ad7
          27352 => x"7c", -- $06ad8
          27353 => x"7c", -- $06ad9
          27354 => x"7c", -- $06ada
          27355 => x"7c", -- $06adb
          27356 => x"7c", -- $06adc
          27357 => x"7c", -- $06add
          27358 => x"7c", -- $06ade
          27359 => x"7c", -- $06adf
          27360 => x"7c", -- $06ae0
          27361 => x"7c", -- $06ae1
          27362 => x"7c", -- $06ae2
          27363 => x"7c", -- $06ae3
          27364 => x"7c", -- $06ae4
          27365 => x"7c", -- $06ae5
          27366 => x"7c", -- $06ae6
          27367 => x"7c", -- $06ae7
          27368 => x"7c", -- $06ae8
          27369 => x"7c", -- $06ae9
          27370 => x"7c", -- $06aea
          27371 => x"7c", -- $06aeb
          27372 => x"7c", -- $06aec
          27373 => x"7c", -- $06aed
          27374 => x"7c", -- $06aee
          27375 => x"7c", -- $06aef
          27376 => x"7c", -- $06af0
          27377 => x"7c", -- $06af1
          27378 => x"7c", -- $06af2
          27379 => x"7c", -- $06af3
          27380 => x"7c", -- $06af4
          27381 => x"7c", -- $06af5
          27382 => x"7c", -- $06af6
          27383 => x"7c", -- $06af7
          27384 => x"7c", -- $06af8
          27385 => x"7c", -- $06af9
          27386 => x"7c", -- $06afa
          27387 => x"7c", -- $06afb
          27388 => x"7c", -- $06afc
          27389 => x"7c", -- $06afd
          27390 => x"7c", -- $06afe
          27391 => x"7c", -- $06aff
          27392 => x"7c", -- $06b00
          27393 => x"7c", -- $06b01
          27394 => x"7c", -- $06b02
          27395 => x"7c", -- $06b03
          27396 => x"7c", -- $06b04
          27397 => x"7c", -- $06b05
          27398 => x"7c", -- $06b06
          27399 => x"7c", -- $06b07
          27400 => x"7c", -- $06b08
          27401 => x"7c", -- $06b09
          27402 => x"7c", -- $06b0a
          27403 => x"7c", -- $06b0b
          27404 => x"7c", -- $06b0c
          27405 => x"7c", -- $06b0d
          27406 => x"7c", -- $06b0e
          27407 => x"7c", -- $06b0f
          27408 => x"7c", -- $06b10
          27409 => x"7c", -- $06b11
          27410 => x"7c", -- $06b12
          27411 => x"7c", -- $06b13
          27412 => x"7c", -- $06b14
          27413 => x"7c", -- $06b15
          27414 => x"7c", -- $06b16
          27415 => x"7c", -- $06b17
          27416 => x"7c", -- $06b18
          27417 => x"7c", -- $06b19
          27418 => x"7c", -- $06b1a
          27419 => x"7c", -- $06b1b
          27420 => x"7c", -- $06b1c
          27421 => x"7c", -- $06b1d
          27422 => x"7c", -- $06b1e
          27423 => x"7c", -- $06b1f
          27424 => x"7c", -- $06b20
          27425 => x"7c", -- $06b21
          27426 => x"7c", -- $06b22
          27427 => x"7c", -- $06b23
          27428 => x"7c", -- $06b24
          27429 => x"7c", -- $06b25
          27430 => x"7c", -- $06b26
          27431 => x"7c", -- $06b27
          27432 => x"7c", -- $06b28
          27433 => x"7c", -- $06b29
          27434 => x"7c", -- $06b2a
          27435 => x"7c", -- $06b2b
          27436 => x"7d", -- $06b2c
          27437 => x"7c", -- $06b2d
          27438 => x"7d", -- $06b2e
          27439 => x"7d", -- $06b2f
          27440 => x"7d", -- $06b30
          27441 => x"7d", -- $06b31
          27442 => x"7d", -- $06b32
          27443 => x"7d", -- $06b33
          27444 => x"7d", -- $06b34
          27445 => x"7d", -- $06b35
          27446 => x"7d", -- $06b36
          27447 => x"7d", -- $06b37
          27448 => x"7d", -- $06b38
          27449 => x"7d", -- $06b39
          27450 => x"7d", -- $06b3a
          27451 => x"7d", -- $06b3b
          27452 => x"7d", -- $06b3c
          27453 => x"7d", -- $06b3d
          27454 => x"7d", -- $06b3e
          27455 => x"7d", -- $06b3f
          27456 => x"7d", -- $06b40
          27457 => x"7d", -- $06b41
          27458 => x"7d", -- $06b42
          27459 => x"7d", -- $06b43
          27460 => x"7d", -- $06b44
          27461 => x"7d", -- $06b45
          27462 => x"7d", -- $06b46
          27463 => x"7d", -- $06b47
          27464 => x"7d", -- $06b48
          27465 => x"7e", -- $06b49
          27466 => x"7e", -- $06b4a
          27467 => x"7e", -- $06b4b
          27468 => x"7e", -- $06b4c
          27469 => x"7e", -- $06b4d
          27470 => x"7e", -- $06b4e
          27471 => x"7e", -- $06b4f
          27472 => x"7e", -- $06b50
          27473 => x"7e", -- $06b51
          27474 => x"7e", -- $06b52
          27475 => x"7e", -- $06b53
          27476 => x"7e", -- $06b54
          27477 => x"7e", -- $06b55
          27478 => x"7e", -- $06b56
          27479 => x"7e", -- $06b57
          27480 => x"7e", -- $06b58
          27481 => x"7e", -- $06b59
          27482 => x"7e", -- $06b5a
          27483 => x"7e", -- $06b5b
          27484 => x"7e", -- $06b5c
          27485 => x"7e", -- $06b5d
          27486 => x"7e", -- $06b5e
          27487 => x"7e", -- $06b5f
          27488 => x"7e", -- $06b60
          27489 => x"7e", -- $06b61
          27490 => x"7f", -- $06b62
          27491 => x"7f", -- $06b63
          27492 => x"7f", -- $06b64
          27493 => x"7f", -- $06b65
          27494 => x"7f", -- $06b66
          27495 => x"7f", -- $06b67
          27496 => x"7f", -- $06b68
          27497 => x"7f", -- $06b69
          27498 => x"7f", -- $06b6a
          27499 => x"7f", -- $06b6b
          27500 => x"7f", -- $06b6c
          27501 => x"7f", -- $06b6d
          27502 => x"7f", -- $06b6e
          27503 => x"7f", -- $06b6f
          27504 => x"7f", -- $06b70
          27505 => x"7f", -- $06b71
          27506 => x"7f", -- $06b72
          27507 => x"7f", -- $06b73
          27508 => x"7f", -- $06b74
          27509 => x"7f", -- $06b75
          27510 => x"7f", -- $06b76
          27511 => x"7f", -- $06b77
          27512 => x"7f", -- $06b78
          27513 => x"7f", -- $06b79
          27514 => x"7f", -- $06b7a
          27515 => x"7f", -- $06b7b
          27516 => x"7f", -- $06b7c
          27517 => x"7f", -- $06b7d
          27518 => x"7f", -- $06b7e
          27519 => x"80", -- $06b7f
          27520 => x"80", -- $06b80
          27521 => x"80", -- $06b81
          27522 => x"7f", -- $06b82
          27523 => x"7f", -- $06b83
          27524 => x"7f", -- $06b84
          27525 => x"80", -- $06b85
          27526 => x"80", -- $06b86
          27527 => x"80", -- $06b87
          27528 => x"80", -- $06b88
          27529 => x"80", -- $06b89
          27530 => x"80", -- $06b8a
          27531 => x"80", -- $06b8b
          27532 => x"80", -- $06b8c
          27533 => x"80", -- $06b8d
          27534 => x"80", -- $06b8e
          27535 => x"80", -- $06b8f
          27536 => x"80", -- $06b90
          27537 => x"80", -- $06b91
          27538 => x"80", -- $06b92
          27539 => x"80", -- $06b93
          27540 => x"80", -- $06b94
          27541 => x"80", -- $06b95
          27542 => x"80", -- $06b96
          27543 => x"80", -- $06b97
          27544 => x"80", -- $06b98
          27545 => x"80", -- $06b99
          27546 => x"80", -- $06b9a
          27547 => x"80", -- $06b9b
          27548 => x"80", -- $06b9c
          27549 => x"80", -- $06b9d
          27550 => x"80", -- $06b9e
          27551 => x"80", -- $06b9f
          27552 => x"80", -- $06ba0
          27553 => x"80", -- $06ba1
          27554 => x"80", -- $06ba2
          27555 => x"80", -- $06ba3
          27556 => x"80", -- $06ba4
          27557 => x"80", -- $06ba5
          27558 => x"80", -- $06ba6
          27559 => x"80", -- $06ba7
          27560 => x"80", -- $06ba8
          27561 => x"80", -- $06ba9
          27562 => x"80", -- $06baa
          27563 => x"80", -- $06bab
          27564 => x"80", -- $06bac
          27565 => x"80", -- $06bad
          27566 => x"80", -- $06bae
          27567 => x"80", -- $06baf
          27568 => x"80", -- $06bb0
          27569 => x"80", -- $06bb1
          27570 => x"80", -- $06bb2
          27571 => x"80", -- $06bb3
          27572 => x"80", -- $06bb4
          27573 => x"81", -- $06bb5
          27574 => x"81", -- $06bb6
          27575 => x"81", -- $06bb7
          27576 => x"81", -- $06bb8
          27577 => x"81", -- $06bb9
          27578 => x"81", -- $06bba
          27579 => x"81", -- $06bbb
          27580 => x"81", -- $06bbc
          27581 => x"81", -- $06bbd
          27582 => x"81", -- $06bbe
          27583 => x"81", -- $06bbf
          27584 => x"81", -- $06bc0
          27585 => x"81", -- $06bc1
          27586 => x"81", -- $06bc2
          27587 => x"81", -- $06bc3
          27588 => x"81", -- $06bc4
          27589 => x"81", -- $06bc5
          27590 => x"81", -- $06bc6
          27591 => x"81", -- $06bc7
          27592 => x"81", -- $06bc8
          27593 => x"81", -- $06bc9
          27594 => x"81", -- $06bca
          27595 => x"81", -- $06bcb
          27596 => x"81", -- $06bcc
          27597 => x"81", -- $06bcd
          27598 => x"81", -- $06bce
          27599 => x"81", -- $06bcf
          27600 => x"81", -- $06bd0
          27601 => x"81", -- $06bd1
          27602 => x"81", -- $06bd2
          27603 => x"81", -- $06bd3
          27604 => x"81", -- $06bd4
          27605 => x"81", -- $06bd5
          27606 => x"81", -- $06bd6
          27607 => x"81", -- $06bd7
          27608 => x"81", -- $06bd8
          27609 => x"81", -- $06bd9
          27610 => x"81", -- $06bda
          27611 => x"82", -- $06bdb
          27612 => x"82", -- $06bdc
          27613 => x"81", -- $06bdd
          27614 => x"81", -- $06bde
          27615 => x"81", -- $06bdf
          27616 => x"81", -- $06be0
          27617 => x"81", -- $06be1
          27618 => x"81", -- $06be2
          27619 => x"81", -- $06be3
          27620 => x"82", -- $06be4
          27621 => x"82", -- $06be5
          27622 => x"82", -- $06be6
          27623 => x"81", -- $06be7
          27624 => x"82", -- $06be8
          27625 => x"82", -- $06be9
          27626 => x"82", -- $06bea
          27627 => x"81", -- $06beb
          27628 => x"81", -- $06bec
          27629 => x"81", -- $06bed
          27630 => x"81", -- $06bee
          27631 => x"81", -- $06bef
          27632 => x"81", -- $06bf0
          27633 => x"81", -- $06bf1
          27634 => x"81", -- $06bf2
          27635 => x"81", -- $06bf3
          27636 => x"81", -- $06bf4
          27637 => x"81", -- $06bf5
          27638 => x"81", -- $06bf6
          27639 => x"81", -- $06bf7
          27640 => x"81", -- $06bf8
          27641 => x"81", -- $06bf9
          27642 => x"81", -- $06bfa
          27643 => x"81", -- $06bfb
          27644 => x"81", -- $06bfc
          27645 => x"81", -- $06bfd
          27646 => x"81", -- $06bfe
          27647 => x"81", -- $06bff
          27648 => x"81", -- $06c00
          27649 => x"81", -- $06c01
          27650 => x"81", -- $06c02
          27651 => x"81", -- $06c03
          27652 => x"81", -- $06c04
          27653 => x"81", -- $06c05
          27654 => x"81", -- $06c06
          27655 => x"81", -- $06c07
          27656 => x"81", -- $06c08
          27657 => x"81", -- $06c09
          27658 => x"81", -- $06c0a
          27659 => x"81", -- $06c0b
          27660 => x"82", -- $06c0c
          27661 => x"82", -- $06c0d
          27662 => x"82", -- $06c0e
          27663 => x"81", -- $06c0f
          27664 => x"81", -- $06c10
          27665 => x"81", -- $06c11
          27666 => x"81", -- $06c12
          27667 => x"81", -- $06c13
          27668 => x"81", -- $06c14
          27669 => x"81", -- $06c15
          27670 => x"81", -- $06c16
          27671 => x"81", -- $06c17
          27672 => x"82", -- $06c18
          27673 => x"82", -- $06c19
          27674 => x"82", -- $06c1a
          27675 => x"82", -- $06c1b
          27676 => x"82", -- $06c1c
          27677 => x"82", -- $06c1d
          27678 => x"82", -- $06c1e
          27679 => x"82", -- $06c1f
          27680 => x"82", -- $06c20
          27681 => x"82", -- $06c21
          27682 => x"82", -- $06c22
          27683 => x"82", -- $06c23
          27684 => x"82", -- $06c24
          27685 => x"82", -- $06c25
          27686 => x"82", -- $06c26
          27687 => x"82", -- $06c27
          27688 => x"82", -- $06c28
          27689 => x"82", -- $06c29
          27690 => x"82", -- $06c2a
          27691 => x"82", -- $06c2b
          27692 => x"82", -- $06c2c
          27693 => x"82", -- $06c2d
          27694 => x"82", -- $06c2e
          27695 => x"82", -- $06c2f
          27696 => x"82", -- $06c30
          27697 => x"82", -- $06c31
          27698 => x"82", -- $06c32
          27699 => x"82", -- $06c33
          27700 => x"82", -- $06c34
          27701 => x"82", -- $06c35
          27702 => x"82", -- $06c36
          27703 => x"82", -- $06c37
          27704 => x"82", -- $06c38
          27705 => x"83", -- $06c39
          27706 => x"82", -- $06c3a
          27707 => x"83", -- $06c3b
          27708 => x"83", -- $06c3c
          27709 => x"83", -- $06c3d
          27710 => x"83", -- $06c3e
          27711 => x"83", -- $06c3f
          27712 => x"83", -- $06c40
          27713 => x"83", -- $06c41
          27714 => x"83", -- $06c42
          27715 => x"83", -- $06c43
          27716 => x"83", -- $06c44
          27717 => x"83", -- $06c45
          27718 => x"83", -- $06c46
          27719 => x"83", -- $06c47
          27720 => x"83", -- $06c48
          27721 => x"83", -- $06c49
          27722 => x"83", -- $06c4a
          27723 => x"83", -- $06c4b
          27724 => x"83", -- $06c4c
          27725 => x"83", -- $06c4d
          27726 => x"83", -- $06c4e
          27727 => x"83", -- $06c4f
          27728 => x"84", -- $06c50
          27729 => x"83", -- $06c51
          27730 => x"83", -- $06c52
          27731 => x"83", -- $06c53
          27732 => x"83", -- $06c54
          27733 => x"84", -- $06c55
          27734 => x"84", -- $06c56
          27735 => x"83", -- $06c57
          27736 => x"84", -- $06c58
          27737 => x"84", -- $06c59
          27738 => x"84", -- $06c5a
          27739 => x"84", -- $06c5b
          27740 => x"84", -- $06c5c
          27741 => x"84", -- $06c5d
          27742 => x"84", -- $06c5e
          27743 => x"84", -- $06c5f
          27744 => x"84", -- $06c60
          27745 => x"84", -- $06c61
          27746 => x"84", -- $06c62
          27747 => x"84", -- $06c63
          27748 => x"84", -- $06c64
          27749 => x"84", -- $06c65
          27750 => x"84", -- $06c66
          27751 => x"84", -- $06c67
          27752 => x"84", -- $06c68
          27753 => x"84", -- $06c69
          27754 => x"84", -- $06c6a
          27755 => x"84", -- $06c6b
          27756 => x"84", -- $06c6c
          27757 => x"84", -- $06c6d
          27758 => x"84", -- $06c6e
          27759 => x"84", -- $06c6f
          27760 => x"84", -- $06c70
          27761 => x"84", -- $06c71
          27762 => x"84", -- $06c72
          27763 => x"84", -- $06c73
          27764 => x"84", -- $06c74
          27765 => x"84", -- $06c75
          27766 => x"84", -- $06c76
          27767 => x"84", -- $06c77
          27768 => x"84", -- $06c78
          27769 => x"84", -- $06c79
          27770 => x"84", -- $06c7a
          27771 => x"84", -- $06c7b
          27772 => x"84", -- $06c7c
          27773 => x"84", -- $06c7d
          27774 => x"84", -- $06c7e
          27775 => x"84", -- $06c7f
          27776 => x"84", -- $06c80
          27777 => x"84", -- $06c81
          27778 => x"84", -- $06c82
          27779 => x"84", -- $06c83
          27780 => x"84", -- $06c84
          27781 => x"84", -- $06c85
          27782 => x"84", -- $06c86
          27783 => x"84", -- $06c87
          27784 => x"84", -- $06c88
          27785 => x"84", -- $06c89
          27786 => x"84", -- $06c8a
          27787 => x"84", -- $06c8b
          27788 => x"84", -- $06c8c
          27789 => x"84", -- $06c8d
          27790 => x"84", -- $06c8e
          27791 => x"84", -- $06c8f
          27792 => x"84", -- $06c90
          27793 => x"84", -- $06c91
          27794 => x"84", -- $06c92
          27795 => x"84", -- $06c93
          27796 => x"84", -- $06c94
          27797 => x"84", -- $06c95
          27798 => x"84", -- $06c96
          27799 => x"84", -- $06c97
          27800 => x"83", -- $06c98
          27801 => x"83", -- $06c99
          27802 => x"83", -- $06c9a
          27803 => x"83", -- $06c9b
          27804 => x"83", -- $06c9c
          27805 => x"83", -- $06c9d
          27806 => x"83", -- $06c9e
          27807 => x"83", -- $06c9f
          27808 => x"83", -- $06ca0
          27809 => x"83", -- $06ca1
          27810 => x"83", -- $06ca2
          27811 => x"83", -- $06ca3
          27812 => x"83", -- $06ca4
          27813 => x"83", -- $06ca5
          27814 => x"83", -- $06ca6
          27815 => x"83", -- $06ca7
          27816 => x"83", -- $06ca8
          27817 => x"83", -- $06ca9
          27818 => x"83", -- $06caa
          27819 => x"83", -- $06cab
          27820 => x"83", -- $06cac
          27821 => x"83", -- $06cad
          27822 => x"83", -- $06cae
          27823 => x"83", -- $06caf
          27824 => x"83", -- $06cb0
          27825 => x"83", -- $06cb1
          27826 => x"83", -- $06cb2
          27827 => x"83", -- $06cb3
          27828 => x"83", -- $06cb4
          27829 => x"83", -- $06cb5
          27830 => x"83", -- $06cb6
          27831 => x"83", -- $06cb7
          27832 => x"83", -- $06cb8
          27833 => x"82", -- $06cb9
          27834 => x"83", -- $06cba
          27835 => x"82", -- $06cbb
          27836 => x"82", -- $06cbc
          27837 => x"82", -- $06cbd
          27838 => x"82", -- $06cbe
          27839 => x"82", -- $06cbf
          27840 => x"82", -- $06cc0
          27841 => x"82", -- $06cc1
          27842 => x"82", -- $06cc2
          27843 => x"82", -- $06cc3
          27844 => x"82", -- $06cc4
          27845 => x"82", -- $06cc5
          27846 => x"82", -- $06cc6
          27847 => x"82", -- $06cc7
          27848 => x"82", -- $06cc8
          27849 => x"82", -- $06cc9
          27850 => x"82", -- $06cca
          27851 => x"82", -- $06ccb
          27852 => x"82", -- $06ccc
          27853 => x"82", -- $06ccd
          27854 => x"82", -- $06cce
          27855 => x"82", -- $06ccf
          27856 => x"82", -- $06cd0
          27857 => x"82", -- $06cd1
          27858 => x"82", -- $06cd2
          27859 => x"82", -- $06cd3
          27860 => x"82", -- $06cd4
          27861 => x"82", -- $06cd5
          27862 => x"82", -- $06cd6
          27863 => x"82", -- $06cd7
          27864 => x"82", -- $06cd8
          27865 => x"82", -- $06cd9
          27866 => x"82", -- $06cda
          27867 => x"82", -- $06cdb
          27868 => x"82", -- $06cdc
          27869 => x"82", -- $06cdd
          27870 => x"82", -- $06cde
          27871 => x"82", -- $06cdf
          27872 => x"82", -- $06ce0
          27873 => x"82", -- $06ce1
          27874 => x"82", -- $06ce2
          27875 => x"82", -- $06ce3
          27876 => x"82", -- $06ce4
          27877 => x"82", -- $06ce5
          27878 => x"82", -- $06ce6
          27879 => x"82", -- $06ce7
          27880 => x"82", -- $06ce8
          27881 => x"82", -- $06ce9
          27882 => x"82", -- $06cea
          27883 => x"82", -- $06ceb
          27884 => x"82", -- $06cec
          27885 => x"82", -- $06ced
          27886 => x"82", -- $06cee
          27887 => x"81", -- $06cef
          27888 => x"81", -- $06cf0
          27889 => x"82", -- $06cf1
          27890 => x"82", -- $06cf2
          27891 => x"81", -- $06cf3
          27892 => x"81", -- $06cf4
          27893 => x"81", -- $06cf5
          27894 => x"81", -- $06cf6
          27895 => x"81", -- $06cf7
          27896 => x"81", -- $06cf8
          27897 => x"81", -- $06cf9
          27898 => x"81", -- $06cfa
          27899 => x"81", -- $06cfb
          27900 => x"81", -- $06cfc
          27901 => x"81", -- $06cfd
          27902 => x"81", -- $06cfe
          27903 => x"81", -- $06cff
          27904 => x"81", -- $06d00
          27905 => x"81", -- $06d01
          27906 => x"81", -- $06d02
          27907 => x"81", -- $06d03
          27908 => x"81", -- $06d04
          27909 => x"81", -- $06d05
          27910 => x"81", -- $06d06
          27911 => x"81", -- $06d07
          27912 => x"81", -- $06d08
          27913 => x"81", -- $06d09
          27914 => x"81", -- $06d0a
          27915 => x"81", -- $06d0b
          27916 => x"81", -- $06d0c
          27917 => x"81", -- $06d0d
          27918 => x"81", -- $06d0e
          27919 => x"81", -- $06d0f
          27920 => x"81", -- $06d10
          27921 => x"81", -- $06d11
          27922 => x"81", -- $06d12
          27923 => x"81", -- $06d13
          27924 => x"81", -- $06d14
          27925 => x"81", -- $06d15
          27926 => x"81", -- $06d16
          27927 => x"81", -- $06d17
          27928 => x"81", -- $06d18
          27929 => x"81", -- $06d19
          27930 => x"80", -- $06d1a
          27931 => x"80", -- $06d1b
          27932 => x"80", -- $06d1c
          27933 => x"81", -- $06d1d
          27934 => x"80", -- $06d1e
          27935 => x"81", -- $06d1f
          27936 => x"81", -- $06d20
          27937 => x"80", -- $06d21
          27938 => x"80", -- $06d22
          27939 => x"80", -- $06d23
          27940 => x"80", -- $06d24
          27941 => x"80", -- $06d25
          27942 => x"80", -- $06d26
          27943 => x"80", -- $06d27
          27944 => x"80", -- $06d28
          27945 => x"80", -- $06d29
          27946 => x"80", -- $06d2a
          27947 => x"80", -- $06d2b
          27948 => x"80", -- $06d2c
          27949 => x"80", -- $06d2d
          27950 => x"80", -- $06d2e
          27951 => x"80", -- $06d2f
          27952 => x"80", -- $06d30
          27953 => x"80", -- $06d31
          27954 => x"80", -- $06d32
          27955 => x"80", -- $06d33
          27956 => x"80", -- $06d34
          27957 => x"80", -- $06d35
          27958 => x"80", -- $06d36
          27959 => x"80", -- $06d37
          27960 => x"80", -- $06d38
          27961 => x"80", -- $06d39
          27962 => x"80", -- $06d3a
          27963 => x"80", -- $06d3b
          27964 => x"80", -- $06d3c
          27965 => x"80", -- $06d3d
          27966 => x"80", -- $06d3e
          27967 => x"80", -- $06d3f
          27968 => x"80", -- $06d40
          27969 => x"80", -- $06d41
          27970 => x"80", -- $06d42
          27971 => x"80", -- $06d43
          27972 => x"80", -- $06d44
          27973 => x"80", -- $06d45
          27974 => x"80", -- $06d46
          27975 => x"80", -- $06d47
          27976 => x"80", -- $06d48
          27977 => x"80", -- $06d49
          27978 => x"80", -- $06d4a
          27979 => x"80", -- $06d4b
          27980 => x"80", -- $06d4c
          27981 => x"80", -- $06d4d
          27982 => x"80", -- $06d4e
          27983 => x"80", -- $06d4f
          27984 => x"80", -- $06d50
          27985 => x"80", -- $06d51
          27986 => x"80", -- $06d52
          27987 => x"80", -- $06d53
          27988 => x"80", -- $06d54
          27989 => x"80", -- $06d55
          27990 => x"80", -- $06d56
          27991 => x"80", -- $06d57
          27992 => x"80", -- $06d58
          27993 => x"80", -- $06d59
          27994 => x"80", -- $06d5a
          27995 => x"80", -- $06d5b
          27996 => x"80", -- $06d5c
          27997 => x"80", -- $06d5d
          27998 => x"80", -- $06d5e
          27999 => x"80", -- $06d5f
          28000 => x"80", -- $06d60
          28001 => x"80", -- $06d61
          28002 => x"80", -- $06d62
          28003 => x"80", -- $06d63
          28004 => x"80", -- $06d64
          28005 => x"80", -- $06d65
          28006 => x"80", -- $06d66
          28007 => x"80", -- $06d67
          28008 => x"80", -- $06d68
          28009 => x"80", -- $06d69
          28010 => x"7f", -- $06d6a
          28011 => x"80", -- $06d6b
          28012 => x"7f", -- $06d6c
          28013 => x"7f", -- $06d6d
          28014 => x"7f", -- $06d6e
          28015 => x"7f", -- $06d6f
          28016 => x"7f", -- $06d70
          28017 => x"7f", -- $06d71
          28018 => x"7f", -- $06d72
          28019 => x"7f", -- $06d73
          28020 => x"7f", -- $06d74
          28021 => x"7f", -- $06d75
          28022 => x"7f", -- $06d76
          28023 => x"7f", -- $06d77
          28024 => x"7f", -- $06d78
          28025 => x"7f", -- $06d79
          28026 => x"7f", -- $06d7a
          28027 => x"7f", -- $06d7b
          28028 => x"7f", -- $06d7c
          28029 => x"7f", -- $06d7d
          28030 => x"7f", -- $06d7e
          28031 => x"7f", -- $06d7f
          28032 => x"7f", -- $06d80
          28033 => x"7f", -- $06d81
          28034 => x"7f", -- $06d82
          28035 => x"7f", -- $06d83
          28036 => x"7f", -- $06d84
          28037 => x"7f", -- $06d85
          28038 => x"7f", -- $06d86
          28039 => x"7f", -- $06d87
          28040 => x"7f", -- $06d88
          28041 => x"7f", -- $06d89
          28042 => x"7f", -- $06d8a
          28043 => x"7f", -- $06d8b
          28044 => x"7f", -- $06d8c
          28045 => x"7f", -- $06d8d
          28046 => x"7f", -- $06d8e
          28047 => x"7e", -- $06d8f
          28048 => x"7e", -- $06d90
          28049 => x"7e", -- $06d91
          28050 => x"7e", -- $06d92
          28051 => x"7e", -- $06d93
          28052 => x"7e", -- $06d94
          28053 => x"7e", -- $06d95
          28054 => x"7e", -- $06d96
          28055 => x"7e", -- $06d97
          28056 => x"7e", -- $06d98
          28057 => x"7e", -- $06d99
          28058 => x"7e", -- $06d9a
          28059 => x"7e", -- $06d9b
          28060 => x"7e", -- $06d9c
          28061 => x"7e", -- $06d9d
          28062 => x"7e", -- $06d9e
          28063 => x"7e", -- $06d9f
          28064 => x"7e", -- $06da0
          28065 => x"7e", -- $06da1
          28066 => x"7e", -- $06da2
          28067 => x"7e", -- $06da3
          28068 => x"7e", -- $06da4
          28069 => x"7e", -- $06da5
          28070 => x"7e", -- $06da6
          28071 => x"7e", -- $06da7
          28072 => x"7e", -- $06da8
          28073 => x"7e", -- $06da9
          28074 => x"7e", -- $06daa
          28075 => x"7e", -- $06dab
          28076 => x"7e", -- $06dac
          28077 => x"7e", -- $06dad
          28078 => x"7e", -- $06dae
          28079 => x"7e", -- $06daf
          28080 => x"7e", -- $06db0
          28081 => x"7e", -- $06db1
          28082 => x"7e", -- $06db2
          28083 => x"7e", -- $06db3
          28084 => x"7e", -- $06db4
          28085 => x"7e", -- $06db5
          28086 => x"7e", -- $06db6
          28087 => x"7e", -- $06db7
          28088 => x"7e", -- $06db8
          28089 => x"7e", -- $06db9
          28090 => x"7e", -- $06dba
          28091 => x"7e", -- $06dbb
          28092 => x"7e", -- $06dbc
          28093 => x"7e", -- $06dbd
          28094 => x"7e", -- $06dbe
          28095 => x"7e", -- $06dbf
          28096 => x"7d", -- $06dc0
          28097 => x"7d", -- $06dc1
          28098 => x"7d", -- $06dc2
          28099 => x"7d", -- $06dc3
          28100 => x"7d", -- $06dc4
          28101 => x"7d", -- $06dc5
          28102 => x"7d", -- $06dc6
          28103 => x"7d", -- $06dc7
          28104 => x"7d", -- $06dc8
          28105 => x"7d", -- $06dc9
          28106 => x"7d", -- $06dca
          28107 => x"7d", -- $06dcb
          28108 => x"7d", -- $06dcc
          28109 => x"7d", -- $06dcd
          28110 => x"7d", -- $06dce
          28111 => x"7d", -- $06dcf
          28112 => x"7d", -- $06dd0
          28113 => x"7d", -- $06dd1
          28114 => x"7d", -- $06dd2
          28115 => x"7d", -- $06dd3
          28116 => x"7d", -- $06dd4
          28117 => x"7d", -- $06dd5
          28118 => x"7d", -- $06dd6
          28119 => x"7d", -- $06dd7
          28120 => x"7d", -- $06dd8
          28121 => x"7d", -- $06dd9
          28122 => x"7d", -- $06dda
          28123 => x"7d", -- $06ddb
          28124 => x"7d", -- $06ddc
          28125 => x"7d", -- $06ddd
          28126 => x"7d", -- $06dde
          28127 => x"7d", -- $06ddf
          28128 => x"7d", -- $06de0
          28129 => x"7d", -- $06de1
          28130 => x"7d", -- $06de2
          28131 => x"7d", -- $06de3
          28132 => x"7d", -- $06de4
          28133 => x"7d", -- $06de5
          28134 => x"7d", -- $06de6
          28135 => x"7d", -- $06de7
          28136 => x"7d", -- $06de8
          28137 => x"7d", -- $06de9
          28138 => x"7d", -- $06dea
          28139 => x"7d", -- $06deb
          28140 => x"7d", -- $06dec
          28141 => x"7d", -- $06ded
          28142 => x"7d", -- $06dee
          28143 => x"7d", -- $06def
          28144 => x"7d", -- $06df0
          28145 => x"7d", -- $06df1
          28146 => x"7d", -- $06df2
          28147 => x"7d", -- $06df3
          28148 => x"7d", -- $06df4
          28149 => x"7d", -- $06df5
          28150 => x"7d", -- $06df6
          28151 => x"7d", -- $06df7
          28152 => x"7d", -- $06df8
          28153 => x"7d", -- $06df9
          28154 => x"7d", -- $06dfa
          28155 => x"7d", -- $06dfb
          28156 => x"7d", -- $06dfc
          28157 => x"7d", -- $06dfd
          28158 => x"7d", -- $06dfe
          28159 => x"7d", -- $06dff
          28160 => x"7d", -- $06e00
          28161 => x"7d", -- $06e01
          28162 => x"7d", -- $06e02
          28163 => x"7d", -- $06e03
          28164 => x"7d", -- $06e04
          28165 => x"7d", -- $06e05
          28166 => x"7d", -- $06e06
          28167 => x"7d", -- $06e07
          28168 => x"7d", -- $06e08
          28169 => x"7d", -- $06e09
          28170 => x"7d", -- $06e0a
          28171 => x"7d", -- $06e0b
          28172 => x"7d", -- $06e0c
          28173 => x"7d", -- $06e0d
          28174 => x"7d", -- $06e0e
          28175 => x"7d", -- $06e0f
          28176 => x"7d", -- $06e10
          28177 => x"7d", -- $06e11
          28178 => x"7d", -- $06e12
          28179 => x"7d", -- $06e13
          28180 => x"7d", -- $06e14
          28181 => x"7d", -- $06e15
          28182 => x"7d", -- $06e16
          28183 => x"7d", -- $06e17
          28184 => x"7d", -- $06e18
          28185 => x"7d", -- $06e19
          28186 => x"7d", -- $06e1a
          28187 => x"7d", -- $06e1b
          28188 => x"7d", -- $06e1c
          28189 => x"7d", -- $06e1d
          28190 => x"7d", -- $06e1e
          28191 => x"7d", -- $06e1f
          28192 => x"7d", -- $06e20
          28193 => x"7d", -- $06e21
          28194 => x"7d", -- $06e22
          28195 => x"7d", -- $06e23
          28196 => x"7d", -- $06e24
          28197 => x"7d", -- $06e25
          28198 => x"7d", -- $06e26
          28199 => x"7d", -- $06e27
          28200 => x"7d", -- $06e28
          28201 => x"7d", -- $06e29
          28202 => x"7d", -- $06e2a
          28203 => x"7d", -- $06e2b
          28204 => x"7d", -- $06e2c
          28205 => x"7d", -- $06e2d
          28206 => x"7d", -- $06e2e
          28207 => x"7d", -- $06e2f
          28208 => x"7d", -- $06e30
          28209 => x"7d", -- $06e31
          28210 => x"7d", -- $06e32
          28211 => x"7d", -- $06e33
          28212 => x"7d", -- $06e34
          28213 => x"7d", -- $06e35
          28214 => x"7d", -- $06e36
          28215 => x"7d", -- $06e37
          28216 => x"7d", -- $06e38
          28217 => x"7d", -- $06e39
          28218 => x"7d", -- $06e3a
          28219 => x"7d", -- $06e3b
          28220 => x"7d", -- $06e3c
          28221 => x"7d", -- $06e3d
          28222 => x"7d", -- $06e3e
          28223 => x"7d", -- $06e3f
          28224 => x"7d", -- $06e40
          28225 => x"7d", -- $06e41
          28226 => x"7d", -- $06e42
          28227 => x"7d", -- $06e43
          28228 => x"7d", -- $06e44
          28229 => x"7d", -- $06e45
          28230 => x"7d", -- $06e46
          28231 => x"7d", -- $06e47
          28232 => x"7d", -- $06e48
          28233 => x"7d", -- $06e49
          28234 => x"7d", -- $06e4a
          28235 => x"7d", -- $06e4b
          28236 => x"7d", -- $06e4c
          28237 => x"7d", -- $06e4d
          28238 => x"7d", -- $06e4e
          28239 => x"7d", -- $06e4f
          28240 => x"7d", -- $06e50
          28241 => x"7d", -- $06e51
          28242 => x"7d", -- $06e52
          28243 => x"7d", -- $06e53
          28244 => x"7d", -- $06e54
          28245 => x"7d", -- $06e55
          28246 => x"7d", -- $06e56
          28247 => x"7d", -- $06e57
          28248 => x"7d", -- $06e58
          28249 => x"7d", -- $06e59
          28250 => x"7d", -- $06e5a
          28251 => x"7d", -- $06e5b
          28252 => x"7d", -- $06e5c
          28253 => x"7d", -- $06e5d
          28254 => x"7d", -- $06e5e
          28255 => x"7d", -- $06e5f
          28256 => x"7d", -- $06e60
          28257 => x"7d", -- $06e61
          28258 => x"7d", -- $06e62
          28259 => x"7d", -- $06e63
          28260 => x"7d", -- $06e64
          28261 => x"7d", -- $06e65
          28262 => x"7d", -- $06e66
          28263 => x"7d", -- $06e67
          28264 => x"7d", -- $06e68
          28265 => x"7d", -- $06e69
          28266 => x"7d", -- $06e6a
          28267 => x"7d", -- $06e6b
          28268 => x"7d", -- $06e6c
          28269 => x"7d", -- $06e6d
          28270 => x"7d", -- $06e6e
          28271 => x"7d", -- $06e6f
          28272 => x"7d", -- $06e70
          28273 => x"7d", -- $06e71
          28274 => x"7e", -- $06e72
          28275 => x"7e", -- $06e73
          28276 => x"7e", -- $06e74
          28277 => x"7e", -- $06e75
          28278 => x"7d", -- $06e76
          28279 => x"7d", -- $06e77
          28280 => x"7d", -- $06e78
          28281 => x"7d", -- $06e79
          28282 => x"7d", -- $06e7a
          28283 => x"7d", -- $06e7b
          28284 => x"7d", -- $06e7c
          28285 => x"7e", -- $06e7d
          28286 => x"7e", -- $06e7e
          28287 => x"7e", -- $06e7f
          28288 => x"7e", -- $06e80
          28289 => x"7e", -- $06e81
          28290 => x"7e", -- $06e82
          28291 => x"7e", -- $06e83
          28292 => x"7e", -- $06e84
          28293 => x"7e", -- $06e85
          28294 => x"7e", -- $06e86
          28295 => x"7e", -- $06e87
          28296 => x"7e", -- $06e88
          28297 => x"7e", -- $06e89
          28298 => x"7e", -- $06e8a
          28299 => x"7e", -- $06e8b
          28300 => x"7e", -- $06e8c
          28301 => x"7e", -- $06e8d
          28302 => x"7e", -- $06e8e
          28303 => x"7e", -- $06e8f
          28304 => x"7e", -- $06e90
          28305 => x"7e", -- $06e91
          28306 => x"7e", -- $06e92
          28307 => x"7e", -- $06e93
          28308 => x"7f", -- $06e94
          28309 => x"7f", -- $06e95
          28310 => x"7f", -- $06e96
          28311 => x"7f", -- $06e97
          28312 => x"7f", -- $06e98
          28313 => x"7f", -- $06e99
          28314 => x"7f", -- $06e9a
          28315 => x"7f", -- $06e9b
          28316 => x"7f", -- $06e9c
          28317 => x"7f", -- $06e9d
          28318 => x"7f", -- $06e9e
          28319 => x"7f", -- $06e9f
          28320 => x"7f", -- $06ea0
          28321 => x"7f", -- $06ea1
          28322 => x"7f", -- $06ea2
          28323 => x"7f", -- $06ea3
          28324 => x"7f", -- $06ea4
          28325 => x"7f", -- $06ea5
          28326 => x"80", -- $06ea6
          28327 => x"80", -- $06ea7
          28328 => x"80", -- $06ea8
          28329 => x"80", -- $06ea9
          28330 => x"80", -- $06eaa
          28331 => x"80", -- $06eab
          28332 => x"80", -- $06eac
          28333 => x"80", -- $06ead
          28334 => x"80", -- $06eae
          28335 => x"80", -- $06eaf
          28336 => x"80", -- $06eb0
          28337 => x"80", -- $06eb1
          28338 => x"80", -- $06eb2
          28339 => x"80", -- $06eb3
          28340 => x"80", -- $06eb4
          28341 => x"80", -- $06eb5
          28342 => x"80", -- $06eb6
          28343 => x"80", -- $06eb7
          28344 => x"80", -- $06eb8
          28345 => x"80", -- $06eb9
          28346 => x"80", -- $06eba
          28347 => x"80", -- $06ebb
          28348 => x"80", -- $06ebc
          28349 => x"80", -- $06ebd
          28350 => x"80", -- $06ebe
          28351 => x"80", -- $06ebf
          28352 => x"80", -- $06ec0
          28353 => x"80", -- $06ec1
          28354 => x"80", -- $06ec2
          28355 => x"80", -- $06ec3
          28356 => x"80", -- $06ec4
          28357 => x"80", -- $06ec5
          28358 => x"80", -- $06ec6
          28359 => x"80", -- $06ec7
          28360 => x"80", -- $06ec8
          28361 => x"80", -- $06ec9
          28362 => x"80", -- $06eca
          28363 => x"80", -- $06ecb
          28364 => x"80", -- $06ecc
          28365 => x"80", -- $06ecd
          28366 => x"80", -- $06ece
          28367 => x"80", -- $06ecf
          28368 => x"81", -- $06ed0
          28369 => x"80", -- $06ed1
          28370 => x"81", -- $06ed2
          28371 => x"81", -- $06ed3
          28372 => x"81", -- $06ed4
          28373 => x"81", -- $06ed5
          28374 => x"81", -- $06ed6
          28375 => x"81", -- $06ed7
          28376 => x"81", -- $06ed8
          28377 => x"81", -- $06ed9
          28378 => x"81", -- $06eda
          28379 => x"81", -- $06edb
          28380 => x"81", -- $06edc
          28381 => x"81", -- $06edd
          28382 => x"81", -- $06ede
          28383 => x"81", -- $06edf
          28384 => x"81", -- $06ee0
          28385 => x"81", -- $06ee1
          28386 => x"81", -- $06ee2
          28387 => x"81", -- $06ee3
          28388 => x"81", -- $06ee4
          28389 => x"81", -- $06ee5
          28390 => x"81", -- $06ee6
          28391 => x"81", -- $06ee7
          28392 => x"82", -- $06ee8
          28393 => x"82", -- $06ee9
          28394 => x"82", -- $06eea
          28395 => x"82", -- $06eeb
          28396 => x"82", -- $06eec
          28397 => x"82", -- $06eed
          28398 => x"82", -- $06eee
          28399 => x"82", -- $06eef
          28400 => x"82", -- $06ef0
          28401 => x"82", -- $06ef1
          28402 => x"82", -- $06ef2
          28403 => x"82", -- $06ef3
          28404 => x"82", -- $06ef4
          28405 => x"82", -- $06ef5
          28406 => x"82", -- $06ef6
          28407 => x"82", -- $06ef7
          28408 => x"82", -- $06ef8
          28409 => x"82", -- $06ef9
          28410 => x"82", -- $06efa
          28411 => x"82", -- $06efb
          28412 => x"82", -- $06efc
          28413 => x"82", -- $06efd
          28414 => x"82", -- $06efe
          28415 => x"82", -- $06eff
          28416 => x"82", -- $06f00
          28417 => x"82", -- $06f01
          28418 => x"82", -- $06f02
          28419 => x"82", -- $06f03
          28420 => x"82", -- $06f04
          28421 => x"82", -- $06f05
          28422 => x"82", -- $06f06
          28423 => x"82", -- $06f07
          28424 => x"82", -- $06f08
          28425 => x"82", -- $06f09
          28426 => x"82", -- $06f0a
          28427 => x"82", -- $06f0b
          28428 => x"82", -- $06f0c
          28429 => x"82", -- $06f0d
          28430 => x"82", -- $06f0e
          28431 => x"82", -- $06f0f
          28432 => x"82", -- $06f10
          28433 => x"82", -- $06f11
          28434 => x"82", -- $06f12
          28435 => x"82", -- $06f13
          28436 => x"82", -- $06f14
          28437 => x"82", -- $06f15
          28438 => x"82", -- $06f16
          28439 => x"82", -- $06f17
          28440 => x"82", -- $06f18
          28441 => x"82", -- $06f19
          28442 => x"82", -- $06f1a
          28443 => x"82", -- $06f1b
          28444 => x"82", -- $06f1c
          28445 => x"82", -- $06f1d
          28446 => x"82", -- $06f1e
          28447 => x"82", -- $06f1f
          28448 => x"82", -- $06f20
          28449 => x"82", -- $06f21
          28450 => x"82", -- $06f22
          28451 => x"82", -- $06f23
          28452 => x"82", -- $06f24
          28453 => x"82", -- $06f25
          28454 => x"82", -- $06f26
          28455 => x"82", -- $06f27
          28456 => x"82", -- $06f28
          28457 => x"82", -- $06f29
          28458 => x"82", -- $06f2a
          28459 => x"82", -- $06f2b
          28460 => x"82", -- $06f2c
          28461 => x"82", -- $06f2d
          28462 => x"82", -- $06f2e
          28463 => x"82", -- $06f2f
          28464 => x"82", -- $06f30
          28465 => x"82", -- $06f31
          28466 => x"82", -- $06f32
          28467 => x"82", -- $06f33
          28468 => x"82", -- $06f34
          28469 => x"82", -- $06f35
          28470 => x"82", -- $06f36
          28471 => x"82", -- $06f37
          28472 => x"82", -- $06f38
          28473 => x"82", -- $06f39
          28474 => x"82", -- $06f3a
          28475 => x"82", -- $06f3b
          28476 => x"82", -- $06f3c
          28477 => x"82", -- $06f3d
          28478 => x"82", -- $06f3e
          28479 => x"82", -- $06f3f
          28480 => x"82", -- $06f40
          28481 => x"82", -- $06f41
          28482 => x"82", -- $06f42
          28483 => x"82", -- $06f43
          28484 => x"82", -- $06f44
          28485 => x"82", -- $06f45
          28486 => x"82", -- $06f46
          28487 => x"82", -- $06f47
          28488 => x"82", -- $06f48
          28489 => x"82", -- $06f49
          28490 => x"82", -- $06f4a
          28491 => x"82", -- $06f4b
          28492 => x"82", -- $06f4c
          28493 => x"82", -- $06f4d
          28494 => x"82", -- $06f4e
          28495 => x"82", -- $06f4f
          28496 => x"82", -- $06f50
          28497 => x"82", -- $06f51
          28498 => x"82", -- $06f52
          28499 => x"82", -- $06f53
          28500 => x"82", -- $06f54
          28501 => x"82", -- $06f55
          28502 => x"82", -- $06f56
          28503 => x"82", -- $06f57
          28504 => x"82", -- $06f58
          28505 => x"82", -- $06f59
          28506 => x"82", -- $06f5a
          28507 => x"82", -- $06f5b
          28508 => x"82", -- $06f5c
          28509 => x"83", -- $06f5d
          28510 => x"83", -- $06f5e
          28511 => x"83", -- $06f5f
          28512 => x"83", -- $06f60
          28513 => x"83", -- $06f61
          28514 => x"83", -- $06f62
          28515 => x"83", -- $06f63
          28516 => x"83", -- $06f64
          28517 => x"83", -- $06f65
          28518 => x"83", -- $06f66
          28519 => x"83", -- $06f67
          28520 => x"83", -- $06f68
          28521 => x"83", -- $06f69
          28522 => x"83", -- $06f6a
          28523 => x"83", -- $06f6b
          28524 => x"83", -- $06f6c
          28525 => x"83", -- $06f6d
          28526 => x"83", -- $06f6e
          28527 => x"83", -- $06f6f
          28528 => x"83", -- $06f70
          28529 => x"83", -- $06f71
          28530 => x"83", -- $06f72
          28531 => x"83", -- $06f73
          28532 => x"83", -- $06f74
          28533 => x"83", -- $06f75
          28534 => x"83", -- $06f76
          28535 => x"83", -- $06f77
          28536 => x"83", -- $06f78
          28537 => x"83", -- $06f79
          28538 => x"83", -- $06f7a
          28539 => x"83", -- $06f7b
          28540 => x"83", -- $06f7c
          28541 => x"83", -- $06f7d
          28542 => x"83", -- $06f7e
          28543 => x"83", -- $06f7f
          28544 => x"83", -- $06f80
          28545 => x"83", -- $06f81
          28546 => x"83", -- $06f82
          28547 => x"83", -- $06f83
          28548 => x"83", -- $06f84
          28549 => x"83", -- $06f85
          28550 => x"83", -- $06f86
          28551 => x"83", -- $06f87
          28552 => x"83", -- $06f88
          28553 => x"83", -- $06f89
          28554 => x"83", -- $06f8a
          28555 => x"83", -- $06f8b
          28556 => x"83", -- $06f8c
          28557 => x"83", -- $06f8d
          28558 => x"83", -- $06f8e
          28559 => x"83", -- $06f8f
          28560 => x"83", -- $06f90
          28561 => x"83", -- $06f91
          28562 => x"83", -- $06f92
          28563 => x"83", -- $06f93
          28564 => x"83", -- $06f94
          28565 => x"83", -- $06f95
          28566 => x"83", -- $06f96
          28567 => x"83", -- $06f97
          28568 => x"83", -- $06f98
          28569 => x"83", -- $06f99
          28570 => x"83", -- $06f9a
          28571 => x"83", -- $06f9b
          28572 => x"83", -- $06f9c
          28573 => x"83", -- $06f9d
          28574 => x"83", -- $06f9e
          28575 => x"83", -- $06f9f
          28576 => x"83", -- $06fa0
          28577 => x"83", -- $06fa1
          28578 => x"83", -- $06fa2
          28579 => x"83", -- $06fa3
          28580 => x"83", -- $06fa4
          28581 => x"83", -- $06fa5
          28582 => x"83", -- $06fa6
          28583 => x"83", -- $06fa7
          28584 => x"83", -- $06fa8
          28585 => x"83", -- $06fa9
          28586 => x"83", -- $06faa
          28587 => x"84", -- $06fab
          28588 => x"83", -- $06fac
          28589 => x"83", -- $06fad
          28590 => x"84", -- $06fae
          28591 => x"83", -- $06faf
          28592 => x"83", -- $06fb0
          28593 => x"83", -- $06fb1
          28594 => x"83", -- $06fb2
          28595 => x"83", -- $06fb3
          28596 => x"83", -- $06fb4
          28597 => x"83", -- $06fb5
          28598 => x"83", -- $06fb6
          28599 => x"83", -- $06fb7
          28600 => x"84", -- $06fb8
          28601 => x"84", -- $06fb9
          28602 => x"83", -- $06fba
          28603 => x"84", -- $06fbb
          28604 => x"84", -- $06fbc
          28605 => x"83", -- $06fbd
          28606 => x"83", -- $06fbe
          28607 => x"83", -- $06fbf
          28608 => x"83", -- $06fc0
          28609 => x"83", -- $06fc1
          28610 => x"83", -- $06fc2
          28611 => x"83", -- $06fc3
          28612 => x"83", -- $06fc4
          28613 => x"83", -- $06fc5
          28614 => x"83", -- $06fc6
          28615 => x"83", -- $06fc7
          28616 => x"83", -- $06fc8
          28617 => x"84", -- $06fc9
          28618 => x"83", -- $06fca
          28619 => x"83", -- $06fcb
          28620 => x"83", -- $06fcc
          28621 => x"83", -- $06fcd
          28622 => x"83", -- $06fce
          28623 => x"83", -- $06fcf
          28624 => x"83", -- $06fd0
          28625 => x"83", -- $06fd1
          28626 => x"83", -- $06fd2
          28627 => x"83", -- $06fd3
          28628 => x"83", -- $06fd4
          28629 => x"83", -- $06fd5
          28630 => x"83", -- $06fd6
          28631 => x"83", -- $06fd7
          28632 => x"83", -- $06fd8
          28633 => x"83", -- $06fd9
          28634 => x"83", -- $06fda
          28635 => x"83", -- $06fdb
          28636 => x"83", -- $06fdc
          28637 => x"83", -- $06fdd
          28638 => x"83", -- $06fde
          28639 => x"83", -- $06fdf
          28640 => x"83", -- $06fe0
          28641 => x"83", -- $06fe1
          28642 => x"83", -- $06fe2
          28643 => x"83", -- $06fe3
          28644 => x"83", -- $06fe4
          28645 => x"83", -- $06fe5
          28646 => x"83", -- $06fe6
          28647 => x"83", -- $06fe7
          28648 => x"83", -- $06fe8
          28649 => x"83", -- $06fe9
          28650 => x"83", -- $06fea
          28651 => x"82", -- $06feb
          28652 => x"82", -- $06fec
          28653 => x"82", -- $06fed
          28654 => x"82", -- $06fee
          28655 => x"82", -- $06fef
          28656 => x"82", -- $06ff0
          28657 => x"82", -- $06ff1
          28658 => x"82", -- $06ff2
          28659 => x"82", -- $06ff3
          28660 => x"82", -- $06ff4
          28661 => x"82", -- $06ff5
          28662 => x"82", -- $06ff6
          28663 => x"82", -- $06ff7
          28664 => x"82", -- $06ff8
          28665 => x"82", -- $06ff9
          28666 => x"82", -- $06ffa
          28667 => x"82", -- $06ffb
          28668 => x"82", -- $06ffc
          28669 => x"82", -- $06ffd
          28670 => x"82", -- $06ffe
          28671 => x"82", -- $06fff
          28672 => x"82", -- $07000
          28673 => x"82", -- $07001
          28674 => x"82", -- $07002
          28675 => x"82", -- $07003
          28676 => x"82", -- $07004
          28677 => x"82", -- $07005
          28678 => x"82", -- $07006
          28679 => x"81", -- $07007
          28680 => x"81", -- $07008
          28681 => x"82", -- $07009
          28682 => x"82", -- $0700a
          28683 => x"81", -- $0700b
          28684 => x"81", -- $0700c
          28685 => x"81", -- $0700d
          28686 => x"81", -- $0700e
          28687 => x"81", -- $0700f
          28688 => x"81", -- $07010
          28689 => x"81", -- $07011
          28690 => x"81", -- $07012
          28691 => x"81", -- $07013
          28692 => x"81", -- $07014
          28693 => x"81", -- $07015
          28694 => x"81", -- $07016
          28695 => x"81", -- $07017
          28696 => x"81", -- $07018
          28697 => x"81", -- $07019
          28698 => x"81", -- $0701a
          28699 => x"81", -- $0701b
          28700 => x"81", -- $0701c
          28701 => x"81", -- $0701d
          28702 => x"81", -- $0701e
          28703 => x"81", -- $0701f
          28704 => x"81", -- $07020
          28705 => x"81", -- $07021
          28706 => x"81", -- $07022
          28707 => x"80", -- $07023
          28708 => x"80", -- $07024
          28709 => x"80", -- $07025
          28710 => x"80", -- $07026
          28711 => x"80", -- $07027
          28712 => x"80", -- $07028
          28713 => x"80", -- $07029
          28714 => x"80", -- $0702a
          28715 => x"80", -- $0702b
          28716 => x"80", -- $0702c
          28717 => x"80", -- $0702d
          28718 => x"80", -- $0702e
          28719 => x"80", -- $0702f
          28720 => x"80", -- $07030
          28721 => x"80", -- $07031
          28722 => x"80", -- $07032
          28723 => x"80", -- $07033
          28724 => x"80", -- $07034
          28725 => x"80", -- $07035
          28726 => x"80", -- $07036
          28727 => x"80", -- $07037
          28728 => x"80", -- $07038
          28729 => x"80", -- $07039
          28730 => x"80", -- $0703a
          28731 => x"80", -- $0703b
          28732 => x"80", -- $0703c
          28733 => x"80", -- $0703d
          28734 => x"80", -- $0703e
          28735 => x"80", -- $0703f
          28736 => x"80", -- $07040
          28737 => x"80", -- $07041
          28738 => x"80", -- $07042
          28739 => x"80", -- $07043
          28740 => x"80", -- $07044
          28741 => x"80", -- $07045
          28742 => x"80", -- $07046
          28743 => x"80", -- $07047
          28744 => x"80", -- $07048
          28745 => x"80", -- $07049
          28746 => x"80", -- $0704a
          28747 => x"80", -- $0704b
          28748 => x"80", -- $0704c
          28749 => x"80", -- $0704d
          28750 => x"80", -- $0704e
          28751 => x"80", -- $0704f
          28752 => x"80", -- $07050
          28753 => x"80", -- $07051
          28754 => x"80", -- $07052
          28755 => x"80", -- $07053
          28756 => x"80", -- $07054
          28757 => x"80", -- $07055
          28758 => x"80", -- $07056
          28759 => x"80", -- $07057
          28760 => x"80", -- $07058
          28761 => x"80", -- $07059
          28762 => x"80", -- $0705a
          28763 => x"80", -- $0705b
          28764 => x"80", -- $0705c
          28765 => x"80", -- $0705d
          28766 => x"80", -- $0705e
          28767 => x"80", -- $0705f
          28768 => x"80", -- $07060
          28769 => x"80", -- $07061
          28770 => x"80", -- $07062
          28771 => x"80", -- $07063
          28772 => x"80", -- $07064
          28773 => x"80", -- $07065
          28774 => x"80", -- $07066
          28775 => x"80", -- $07067
          28776 => x"80", -- $07068
          28777 => x"80", -- $07069
          28778 => x"80", -- $0706a
          28779 => x"80", -- $0706b
          28780 => x"80", -- $0706c
          28781 => x"80", -- $0706d
          28782 => x"80", -- $0706e
          28783 => x"80", -- $0706f
          28784 => x"80", -- $07070
          28785 => x"80", -- $07071
          28786 => x"80", -- $07072
          28787 => x"80", -- $07073
          28788 => x"80", -- $07074
          28789 => x"80", -- $07075
          28790 => x"80", -- $07076
          28791 => x"80", -- $07077
          28792 => x"80", -- $07078
          28793 => x"80", -- $07079
          28794 => x"80", -- $0707a
          28795 => x"80", -- $0707b
          28796 => x"80", -- $0707c
          28797 => x"80", -- $0707d
          28798 => x"80", -- $0707e
          28799 => x"80", -- $0707f
          28800 => x"80", -- $07080
          28801 => x"80", -- $07081
          28802 => x"80", -- $07082
          28803 => x"80", -- $07083
          28804 => x"80", -- $07084
          28805 => x"7f", -- $07085
          28806 => x"7f", -- $07086
          28807 => x"80", -- $07087
          28808 => x"80", -- $07088
          28809 => x"80", -- $07089
          28810 => x"80", -- $0708a
          28811 => x"80", -- $0708b
          28812 => x"80", -- $0708c
          28813 => x"80", -- $0708d
          28814 => x"7f", -- $0708e
          28815 => x"7f", -- $0708f
          28816 => x"7f", -- $07090
          28817 => x"7f", -- $07091
          28818 => x"7f", -- $07092
          28819 => x"7f", -- $07093
          28820 => x"7f", -- $07094
          28821 => x"7f", -- $07095
          28822 => x"7f", -- $07096
          28823 => x"7f", -- $07097
          28824 => x"7f", -- $07098
          28825 => x"7f", -- $07099
          28826 => x"7f", -- $0709a
          28827 => x"7f", -- $0709b
          28828 => x"7f", -- $0709c
          28829 => x"7f", -- $0709d
          28830 => x"7f", -- $0709e
          28831 => x"7f", -- $0709f
          28832 => x"7f", -- $070a0
          28833 => x"7f", -- $070a1
          28834 => x"7f", -- $070a2
          28835 => x"7f", -- $070a3
          28836 => x"7f", -- $070a4
          28837 => x"7f", -- $070a5
          28838 => x"7f", -- $070a6
          28839 => x"7f", -- $070a7
          28840 => x"7f", -- $070a8
          28841 => x"7f", -- $070a9
          28842 => x"7f", -- $070aa
          28843 => x"7f", -- $070ab
          28844 => x"7f", -- $070ac
          28845 => x"7f", -- $070ad
          28846 => x"7f", -- $070ae
          28847 => x"7f", -- $070af
          28848 => x"7f", -- $070b0
          28849 => x"7f", -- $070b1
          28850 => x"7f", -- $070b2
          28851 => x"7f", -- $070b3
          28852 => x"7f", -- $070b4
          28853 => x"7f", -- $070b5
          28854 => x"7f", -- $070b6
          28855 => x"7f", -- $070b7
          28856 => x"7e", -- $070b8
          28857 => x"7e", -- $070b9
          28858 => x"7e", -- $070ba
          28859 => x"7f", -- $070bb
          28860 => x"7f", -- $070bc
          28861 => x"7f", -- $070bd
          28862 => x"7e", -- $070be
          28863 => x"7e", -- $070bf
          28864 => x"7f", -- $070c0
          28865 => x"7e", -- $070c1
          28866 => x"7e", -- $070c2
          28867 => x"7e", -- $070c3
          28868 => x"7e", -- $070c4
          28869 => x"7e", -- $070c5
          28870 => x"7e", -- $070c6
          28871 => x"7e", -- $070c7
          28872 => x"7e", -- $070c8
          28873 => x"7e", -- $070c9
          28874 => x"7e", -- $070ca
          28875 => x"7e", -- $070cb
          28876 => x"7e", -- $070cc
          28877 => x"7e", -- $070cd
          28878 => x"7e", -- $070ce
          28879 => x"7e", -- $070cf
          28880 => x"7e", -- $070d0
          28881 => x"7e", -- $070d1
          28882 => x"7e", -- $070d2
          28883 => x"7e", -- $070d3
          28884 => x"7e", -- $070d4
          28885 => x"7d", -- $070d5
          28886 => x"7e", -- $070d6
          28887 => x"7e", -- $070d7
          28888 => x"7e", -- $070d8
          28889 => x"7e", -- $070d9
          28890 => x"7e", -- $070da
          28891 => x"7d", -- $070db
          28892 => x"7d", -- $070dc
          28893 => x"7d", -- $070dd
          28894 => x"7d", -- $070de
          28895 => x"7d", -- $070df
          28896 => x"7d", -- $070e0
          28897 => x"7d", -- $070e1
          28898 => x"7d", -- $070e2
          28899 => x"7d", -- $070e3
          28900 => x"7d", -- $070e4
          28901 => x"7d", -- $070e5
          28902 => x"7d", -- $070e6
          28903 => x"7d", -- $070e7
          28904 => x"7d", -- $070e8
          28905 => x"7d", -- $070e9
          28906 => x"7d", -- $070ea
          28907 => x"7d", -- $070eb
          28908 => x"7d", -- $070ec
          28909 => x"7d", -- $070ed
          28910 => x"7d", -- $070ee
          28911 => x"7d", -- $070ef
          28912 => x"7d", -- $070f0
          28913 => x"7d", -- $070f1
          28914 => x"7d", -- $070f2
          28915 => x"7d", -- $070f3
          28916 => x"7d", -- $070f4
          28917 => x"7c", -- $070f5
          28918 => x"7d", -- $070f6
          28919 => x"7c", -- $070f7
          28920 => x"7c", -- $070f8
          28921 => x"7c", -- $070f9
          28922 => x"7c", -- $070fa
          28923 => x"7c", -- $070fb
          28924 => x"7c", -- $070fc
          28925 => x"7c", -- $070fd
          28926 => x"7c", -- $070fe
          28927 => x"7c", -- $070ff
          28928 => x"7c", -- $07100
          28929 => x"7c", -- $07101
          28930 => x"7c", -- $07102
          28931 => x"7c", -- $07103
          28932 => x"7c", -- $07104
          28933 => x"7c", -- $07105
          28934 => x"7c", -- $07106
          28935 => x"7c", -- $07107
          28936 => x"7c", -- $07108
          28937 => x"7c", -- $07109
          28938 => x"7c", -- $0710a
          28939 => x"7c", -- $0710b
          28940 => x"7c", -- $0710c
          28941 => x"7c", -- $0710d
          28942 => x"7c", -- $0710e
          28943 => x"7c", -- $0710f
          28944 => x"7c", -- $07110
          28945 => x"7c", -- $07111
          28946 => x"7c", -- $07112
          28947 => x"7c", -- $07113
          28948 => x"7c", -- $07114
          28949 => x"7c", -- $07115
          28950 => x"7c", -- $07116
          28951 => x"7c", -- $07117
          28952 => x"7c", -- $07118
          28953 => x"7c", -- $07119
          28954 => x"7c", -- $0711a
          28955 => x"7c", -- $0711b
          28956 => x"7c", -- $0711c
          28957 => x"7c", -- $0711d
          28958 => x"7c", -- $0711e
          28959 => x"7c", -- $0711f
          28960 => x"7c", -- $07120
          28961 => x"7c", -- $07121
          28962 => x"7c", -- $07122
          28963 => x"7c", -- $07123
          28964 => x"7c", -- $07124
          28965 => x"7c", -- $07125
          28966 => x"7c", -- $07126
          28967 => x"7c", -- $07127
          28968 => x"7c", -- $07128
          28969 => x"7c", -- $07129
          28970 => x"7c", -- $0712a
          28971 => x"7c", -- $0712b
          28972 => x"7c", -- $0712c
          28973 => x"7c", -- $0712d
          28974 => x"7c", -- $0712e
          28975 => x"7c", -- $0712f
          28976 => x"7c", -- $07130
          28977 => x"7c", -- $07131
          28978 => x"7c", -- $07132
          28979 => x"7c", -- $07133
          28980 => x"7c", -- $07134
          28981 => x"7c", -- $07135
          28982 => x"7c", -- $07136
          28983 => x"7c", -- $07137
          28984 => x"7c", -- $07138
          28985 => x"7c", -- $07139
          28986 => x"7c", -- $0713a
          28987 => x"7c", -- $0713b
          28988 => x"7c", -- $0713c
          28989 => x"7c", -- $0713d
          28990 => x"7d", -- $0713e
          28991 => x"7d", -- $0713f
          28992 => x"7d", -- $07140
          28993 => x"7d", -- $07141
          28994 => x"7d", -- $07142
          28995 => x"7d", -- $07143
          28996 => x"7d", -- $07144
          28997 => x"7d", -- $07145
          28998 => x"7d", -- $07146
          28999 => x"7d", -- $07147
          29000 => x"7d", -- $07148
          29001 => x"7d", -- $07149
          29002 => x"7d", -- $0714a
          29003 => x"7d", -- $0714b
          29004 => x"7d", -- $0714c
          29005 => x"7d", -- $0714d
          29006 => x"7d", -- $0714e
          29007 => x"7d", -- $0714f
          29008 => x"7d", -- $07150
          29009 => x"7d", -- $07151
          29010 => x"7d", -- $07152
          29011 => x"7d", -- $07153
          29012 => x"7d", -- $07154
          29013 => x"7d", -- $07155
          29014 => x"7d", -- $07156
          29015 => x"7d", -- $07157
          29016 => x"7d", -- $07158
          29017 => x"7d", -- $07159
          29018 => x"7d", -- $0715a
          29019 => x"7d", -- $0715b
          29020 => x"7d", -- $0715c
          29021 => x"7d", -- $0715d
          29022 => x"7d", -- $0715e
          29023 => x"7d", -- $0715f
          29024 => x"7d", -- $07160
          29025 => x"7d", -- $07161
          29026 => x"7d", -- $07162
          29027 => x"7d", -- $07163
          29028 => x"7d", -- $07164
          29029 => x"7d", -- $07165
          29030 => x"7d", -- $07166
          29031 => x"7e", -- $07167
          29032 => x"7e", -- $07168
          29033 => x"7e", -- $07169
          29034 => x"7e", -- $0716a
          29035 => x"7e", -- $0716b
          29036 => x"7e", -- $0716c
          29037 => x"7e", -- $0716d
          29038 => x"7e", -- $0716e
          29039 => x"7e", -- $0716f
          29040 => x"7e", -- $07170
          29041 => x"7e", -- $07171
          29042 => x"7e", -- $07172
          29043 => x"7e", -- $07173
          29044 => x"7e", -- $07174
          29045 => x"7e", -- $07175
          29046 => x"7e", -- $07176
          29047 => x"7e", -- $07177
          29048 => x"7e", -- $07178
          29049 => x"7e", -- $07179
          29050 => x"7e", -- $0717a
          29051 => x"7e", -- $0717b
          29052 => x"7e", -- $0717c
          29053 => x"7e", -- $0717d
          29054 => x"7e", -- $0717e
          29055 => x"7e", -- $0717f
          29056 => x"7e", -- $07180
          29057 => x"7e", -- $07181
          29058 => x"7e", -- $07182
          29059 => x"7e", -- $07183
          29060 => x"7e", -- $07184
          29061 => x"7e", -- $07185
          29062 => x"7e", -- $07186
          29063 => x"7e", -- $07187
          29064 => x"7e", -- $07188
          29065 => x"7e", -- $07189
          29066 => x"7e", -- $0718a
          29067 => x"7e", -- $0718b
          29068 => x"7e", -- $0718c
          29069 => x"7e", -- $0718d
          29070 => x"7e", -- $0718e
          29071 => x"7e", -- $0718f
          29072 => x"7e", -- $07190
          29073 => x"7f", -- $07191
          29074 => x"7e", -- $07192
          29075 => x"7e", -- $07193
          29076 => x"7e", -- $07194
          29077 => x"7e", -- $07195
          29078 => x"7e", -- $07196
          29079 => x"7e", -- $07197
          29080 => x"7e", -- $07198
          29081 => x"7e", -- $07199
          29082 => x"7f", -- $0719a
          29083 => x"7e", -- $0719b
          29084 => x"7e", -- $0719c
          29085 => x"7e", -- $0719d
          29086 => x"7f", -- $0719e
          29087 => x"7f", -- $0719f
          29088 => x"7f", -- $071a0
          29089 => x"7e", -- $071a1
          29090 => x"7e", -- $071a2
          29091 => x"7f", -- $071a3
          29092 => x"7e", -- $071a4
          29093 => x"7e", -- $071a5
          29094 => x"7e", -- $071a6
          29095 => x"7f", -- $071a7
          29096 => x"7f", -- $071a8
          29097 => x"7e", -- $071a9
          29098 => x"7f", -- $071aa
          29099 => x"7f", -- $071ab
          29100 => x"7f", -- $071ac
          29101 => x"7f", -- $071ad
          29102 => x"7f", -- $071ae
          29103 => x"7f", -- $071af
          29104 => x"7f", -- $071b0
          29105 => x"7f", -- $071b1
          29106 => x"7f", -- $071b2
          29107 => x"7f", -- $071b3
          29108 => x"7f", -- $071b4
          29109 => x"7f", -- $071b5
          29110 => x"7f", -- $071b6
          29111 => x"7f", -- $071b7
          29112 => x"7f", -- $071b8
          29113 => x"7f", -- $071b9
          29114 => x"7f", -- $071ba
          29115 => x"7f", -- $071bb
          29116 => x"7f", -- $071bc
          29117 => x"7f", -- $071bd
          29118 => x"7f", -- $071be
          29119 => x"7f", -- $071bf
          29120 => x"7f", -- $071c0
          29121 => x"7f", -- $071c1
          29122 => x"7f", -- $071c2
          29123 => x"7f", -- $071c3
          29124 => x"7f", -- $071c4
          29125 => x"7f", -- $071c5
          29126 => x"7f", -- $071c6
          29127 => x"7f", -- $071c7
          29128 => x"80", -- $071c8
          29129 => x"80", -- $071c9
          29130 => x"80", -- $071ca
          29131 => x"80", -- $071cb
          29132 => x"80", -- $071cc
          29133 => x"80", -- $071cd
          29134 => x"80", -- $071ce
          29135 => x"80", -- $071cf
          29136 => x"80", -- $071d0
          29137 => x"80", -- $071d1
          29138 => x"80", -- $071d2
          29139 => x"80", -- $071d3
          29140 => x"80", -- $071d4
          29141 => x"80", -- $071d5
          29142 => x"80", -- $071d6
          29143 => x"80", -- $071d7
          29144 => x"80", -- $071d8
          29145 => x"80", -- $071d9
          29146 => x"80", -- $071da
          29147 => x"80", -- $071db
          29148 => x"80", -- $071dc
          29149 => x"80", -- $071dd
          29150 => x"80", -- $071de
          29151 => x"80", -- $071df
          29152 => x"80", -- $071e0
          29153 => x"80", -- $071e1
          29154 => x"80", -- $071e2
          29155 => x"80", -- $071e3
          29156 => x"80", -- $071e4
          29157 => x"80", -- $071e5
          29158 => x"80", -- $071e6
          29159 => x"80", -- $071e7
          29160 => x"80", -- $071e8
          29161 => x"80", -- $071e9
          29162 => x"80", -- $071ea
          29163 => x"80", -- $071eb
          29164 => x"80", -- $071ec
          29165 => x"80", -- $071ed
          29166 => x"80", -- $071ee
          29167 => x"80", -- $071ef
          29168 => x"80", -- $071f0
          29169 => x"80", -- $071f1
          29170 => x"80", -- $071f2
          29171 => x"80", -- $071f3
          29172 => x"80", -- $071f4
          29173 => x"80", -- $071f5
          29174 => x"80", -- $071f6
          29175 => x"80", -- $071f7
          29176 => x"80", -- $071f8
          29177 => x"80", -- $071f9
          29178 => x"80", -- $071fa
          29179 => x"80", -- $071fb
          29180 => x"80", -- $071fc
          29181 => x"80", -- $071fd
          29182 => x"80", -- $071fe
          29183 => x"80", -- $071ff
          29184 => x"80", -- $07200
          29185 => x"80", -- $07201
          29186 => x"81", -- $07202
          29187 => x"81", -- $07203
          29188 => x"81", -- $07204
          29189 => x"81", -- $07205
          29190 => x"81", -- $07206
          29191 => x"81", -- $07207
          29192 => x"81", -- $07208
          29193 => x"81", -- $07209
          29194 => x"81", -- $0720a
          29195 => x"81", -- $0720b
          29196 => x"81", -- $0720c
          29197 => x"81", -- $0720d
          29198 => x"81", -- $0720e
          29199 => x"81", -- $0720f
          29200 => x"81", -- $07210
          29201 => x"81", -- $07211
          29202 => x"81", -- $07212
          29203 => x"81", -- $07213
          29204 => x"81", -- $07214
          29205 => x"81", -- $07215
          29206 => x"81", -- $07216
          29207 => x"81", -- $07217
          29208 => x"81", -- $07218
          29209 => x"81", -- $07219
          29210 => x"81", -- $0721a
          29211 => x"81", -- $0721b
          29212 => x"81", -- $0721c
          29213 => x"82", -- $0721d
          29214 => x"81", -- $0721e
          29215 => x"82", -- $0721f
          29216 => x"82", -- $07220
          29217 => x"81", -- $07221
          29218 => x"81", -- $07222
          29219 => x"82", -- $07223
          29220 => x"82", -- $07224
          29221 => x"82", -- $07225
          29222 => x"82", -- $07226
          29223 => x"82", -- $07227
          29224 => x"82", -- $07228
          29225 => x"82", -- $07229
          29226 => x"82", -- $0722a
          29227 => x"82", -- $0722b
          29228 => x"82", -- $0722c
          29229 => x"82", -- $0722d
          29230 => x"82", -- $0722e
          29231 => x"82", -- $0722f
          29232 => x"82", -- $07230
          29233 => x"82", -- $07231
          29234 => x"82", -- $07232
          29235 => x"82", -- $07233
          29236 => x"82", -- $07234
          29237 => x"82", -- $07235
          29238 => x"82", -- $07236
          29239 => x"82", -- $07237
          29240 => x"82", -- $07238
          29241 => x"82", -- $07239
          29242 => x"82", -- $0723a
          29243 => x"82", -- $0723b
          29244 => x"82", -- $0723c
          29245 => x"82", -- $0723d
          29246 => x"82", -- $0723e
          29247 => x"82", -- $0723f
          29248 => x"82", -- $07240
          29249 => x"82", -- $07241
          29250 => x"82", -- $07242
          29251 => x"82", -- $07243
          29252 => x"82", -- $07244
          29253 => x"82", -- $07245
          29254 => x"82", -- $07246
          29255 => x"83", -- $07247
          29256 => x"82", -- $07248
          29257 => x"83", -- $07249
          29258 => x"82", -- $0724a
          29259 => x"83", -- $0724b
          29260 => x"83", -- $0724c
          29261 => x"83", -- $0724d
          29262 => x"83", -- $0724e
          29263 => x"83", -- $0724f
          29264 => x"83", -- $07250
          29265 => x"83", -- $07251
          29266 => x"83", -- $07252
          29267 => x"83", -- $07253
          29268 => x"83", -- $07254
          29269 => x"83", -- $07255
          29270 => x"83", -- $07256
          29271 => x"83", -- $07257
          29272 => x"83", -- $07258
          29273 => x"83", -- $07259
          29274 => x"83", -- $0725a
          29275 => x"83", -- $0725b
          29276 => x"83", -- $0725c
          29277 => x"83", -- $0725d
          29278 => x"83", -- $0725e
          29279 => x"83", -- $0725f
          29280 => x"83", -- $07260
          29281 => x"83", -- $07261
          29282 => x"83", -- $07262
          29283 => x"83", -- $07263
          29284 => x"83", -- $07264
          29285 => x"83", -- $07265
          29286 => x"83", -- $07266
          29287 => x"83", -- $07267
          29288 => x"83", -- $07268
          29289 => x"83", -- $07269
          29290 => x"83", -- $0726a
          29291 => x"83", -- $0726b
          29292 => x"83", -- $0726c
          29293 => x"83", -- $0726d
          29294 => x"83", -- $0726e
          29295 => x"83", -- $0726f
          29296 => x"83", -- $07270
          29297 => x"83", -- $07271
          29298 => x"83", -- $07272
          29299 => x"83", -- $07273
          29300 => x"83", -- $07274
          29301 => x"83", -- $07275
          29302 => x"83", -- $07276
          29303 => x"83", -- $07277
          29304 => x"83", -- $07278
          29305 => x"84", -- $07279
          29306 => x"84", -- $0727a
          29307 => x"84", -- $0727b
          29308 => x"84", -- $0727c
          29309 => x"84", -- $0727d
          29310 => x"84", -- $0727e
          29311 => x"84", -- $0727f
          29312 => x"83", -- $07280
          29313 => x"83", -- $07281
          29314 => x"84", -- $07282
          29315 => x"83", -- $07283
          29316 => x"84", -- $07284
          29317 => x"84", -- $07285
          29318 => x"84", -- $07286
          29319 => x"84", -- $07287
          29320 => x"84", -- $07288
          29321 => x"84", -- $07289
          29322 => x"84", -- $0728a
          29323 => x"84", -- $0728b
          29324 => x"83", -- $0728c
          29325 => x"83", -- $0728d
          29326 => x"83", -- $0728e
          29327 => x"83", -- $0728f
          29328 => x"83", -- $07290
          29329 => x"83", -- $07291
          29330 => x"83", -- $07292
          29331 => x"83", -- $07293
          29332 => x"83", -- $07294
          29333 => x"84", -- $07295
          29334 => x"84", -- $07296
          29335 => x"84", -- $07297
          29336 => x"84", -- $07298
          29337 => x"83", -- $07299
          29338 => x"83", -- $0729a
          29339 => x"83", -- $0729b
          29340 => x"83", -- $0729c
          29341 => x"83", -- $0729d
          29342 => x"83", -- $0729e
          29343 => x"83", -- $0729f
          29344 => x"84", -- $072a0
          29345 => x"84", -- $072a1
          29346 => x"84", -- $072a2
          29347 => x"84", -- $072a3
          29348 => x"83", -- $072a4
          29349 => x"83", -- $072a5
          29350 => x"83", -- $072a6
          29351 => x"83", -- $072a7
          29352 => x"83", -- $072a8
          29353 => x"83", -- $072a9
          29354 => x"83", -- $072aa
          29355 => x"83", -- $072ab
          29356 => x"83", -- $072ac
          29357 => x"83", -- $072ad
          29358 => x"83", -- $072ae
          29359 => x"83", -- $072af
          29360 => x"83", -- $072b0
          29361 => x"83", -- $072b1
          29362 => x"83", -- $072b2
          29363 => x"83", -- $072b3
          29364 => x"83", -- $072b4
          29365 => x"83", -- $072b5
          29366 => x"83", -- $072b6
          29367 => x"83", -- $072b7
          29368 => x"83", -- $072b8
          29369 => x"83", -- $072b9
          29370 => x"83", -- $072ba
          29371 => x"83", -- $072bb
          29372 => x"83", -- $072bc
          29373 => x"83", -- $072bd
          29374 => x"83", -- $072be
          29375 => x"83", -- $072bf
          29376 => x"83", -- $072c0
          29377 => x"83", -- $072c1
          29378 => x"83", -- $072c2
          29379 => x"83", -- $072c3
          29380 => x"83", -- $072c4
          29381 => x"83", -- $072c5
          29382 => x"83", -- $072c6
          29383 => x"83", -- $072c7
          29384 => x"83", -- $072c8
          29385 => x"83", -- $072c9
          29386 => x"83", -- $072ca
          29387 => x"83", -- $072cb
          29388 => x"83", -- $072cc
          29389 => x"83", -- $072cd
          29390 => x"83", -- $072ce
          29391 => x"83", -- $072cf
          29392 => x"83", -- $072d0
          29393 => x"83", -- $072d1
          29394 => x"83", -- $072d2
          29395 => x"83", -- $072d3
          29396 => x"83", -- $072d4
          29397 => x"83", -- $072d5
          29398 => x"83", -- $072d6
          29399 => x"83", -- $072d7
          29400 => x"83", -- $072d8
          29401 => x"83", -- $072d9
          29402 => x"83", -- $072da
          29403 => x"83", -- $072db
          29404 => x"83", -- $072dc
          29405 => x"83", -- $072dd
          29406 => x"83", -- $072de
          29407 => x"83", -- $072df
          29408 => x"83", -- $072e0
          29409 => x"83", -- $072e1
          29410 => x"83", -- $072e2
          29411 => x"83", -- $072e3
          29412 => x"83", -- $072e4
          29413 => x"83", -- $072e5
          29414 => x"83", -- $072e6
          29415 => x"83", -- $072e7
          29416 => x"83", -- $072e8
          29417 => x"83", -- $072e9
          29418 => x"83", -- $072ea
          29419 => x"83", -- $072eb
          29420 => x"83", -- $072ec
          29421 => x"82", -- $072ed
          29422 => x"82", -- $072ee
          29423 => x"83", -- $072ef
          29424 => x"83", -- $072f0
          29425 => x"82", -- $072f1
          29426 => x"82", -- $072f2
          29427 => x"82", -- $072f3
          29428 => x"82", -- $072f4
          29429 => x"82", -- $072f5
          29430 => x"82", -- $072f6
          29431 => x"82", -- $072f7
          29432 => x"82", -- $072f8
          29433 => x"82", -- $072f9
          29434 => x"82", -- $072fa
          29435 => x"82", -- $072fb
          29436 => x"82", -- $072fc
          29437 => x"83", -- $072fd
          29438 => x"82", -- $072fe
          29439 => x"83", -- $072ff
          29440 => x"83", -- $07300
          29441 => x"83", -- $07301
          29442 => x"83", -- $07302
          29443 => x"82", -- $07303
          29444 => x"82", -- $07304
          29445 => x"83", -- $07305
          29446 => x"83", -- $07306
          29447 => x"83", -- $07307
          29448 => x"83", -- $07308
          29449 => x"83", -- $07309
          29450 => x"83", -- $0730a
          29451 => x"82", -- $0730b
          29452 => x"82", -- $0730c
          29453 => x"82", -- $0730d
          29454 => x"82", -- $0730e
          29455 => x"82", -- $0730f
          29456 => x"82", -- $07310
          29457 => x"82", -- $07311
          29458 => x"82", -- $07312
          29459 => x"82", -- $07313
          29460 => x"82", -- $07314
          29461 => x"82", -- $07315
          29462 => x"82", -- $07316
          29463 => x"82", -- $07317
          29464 => x"82", -- $07318
          29465 => x"82", -- $07319
          29466 => x"82", -- $0731a
          29467 => x"82", -- $0731b
          29468 => x"82", -- $0731c
          29469 => x"82", -- $0731d
          29470 => x"82", -- $0731e
          29471 => x"82", -- $0731f
          29472 => x"82", -- $07320
          29473 => x"82", -- $07321
          29474 => x"82", -- $07322
          29475 => x"82", -- $07323
          29476 => x"82", -- $07324
          29477 => x"82", -- $07325
          29478 => x"82", -- $07326
          29479 => x"82", -- $07327
          29480 => x"82", -- $07328
          29481 => x"82", -- $07329
          29482 => x"82", -- $0732a
          29483 => x"82", -- $0732b
          29484 => x"82", -- $0732c
          29485 => x"82", -- $0732d
          29486 => x"81", -- $0732e
          29487 => x"81", -- $0732f
          29488 => x"82", -- $07330
          29489 => x"82", -- $07331
          29490 => x"81", -- $07332
          29491 => x"81", -- $07333
          29492 => x"82", -- $07334
          29493 => x"81", -- $07335
          29494 => x"81", -- $07336
          29495 => x"81", -- $07337
          29496 => x"81", -- $07338
          29497 => x"81", -- $07339
          29498 => x"81", -- $0733a
          29499 => x"81", -- $0733b
          29500 => x"81", -- $0733c
          29501 => x"81", -- $0733d
          29502 => x"81", -- $0733e
          29503 => x"81", -- $0733f
          29504 => x"81", -- $07340
          29505 => x"81", -- $07341
          29506 => x"81", -- $07342
          29507 => x"81", -- $07343
          29508 => x"81", -- $07344
          29509 => x"81", -- $07345
          29510 => x"81", -- $07346
          29511 => x"80", -- $07347
          29512 => x"81", -- $07348
          29513 => x"80", -- $07349
          29514 => x"80", -- $0734a
          29515 => x"80", -- $0734b
          29516 => x"80", -- $0734c
          29517 => x"80", -- $0734d
          29518 => x"80", -- $0734e
          29519 => x"80", -- $0734f
          29520 => x"80", -- $07350
          29521 => x"80", -- $07351
          29522 => x"80", -- $07352
          29523 => x"80", -- $07353
          29524 => x"80", -- $07354
          29525 => x"80", -- $07355
          29526 => x"80", -- $07356
          29527 => x"80", -- $07357
          29528 => x"80", -- $07358
          29529 => x"80", -- $07359
          29530 => x"80", -- $0735a
          29531 => x"80", -- $0735b
          29532 => x"80", -- $0735c
          29533 => x"80", -- $0735d
          29534 => x"80", -- $0735e
          29535 => x"80", -- $0735f
          29536 => x"80", -- $07360
          29537 => x"80", -- $07361
          29538 => x"80", -- $07362
          29539 => x"80", -- $07363
          29540 => x"80", -- $07364
          29541 => x"80", -- $07365
          29542 => x"80", -- $07366
          29543 => x"80", -- $07367
          29544 => x"80", -- $07368
          29545 => x"80", -- $07369
          29546 => x"80", -- $0736a
          29547 => x"80", -- $0736b
          29548 => x"80", -- $0736c
          29549 => x"80", -- $0736d
          29550 => x"80", -- $0736e
          29551 => x"80", -- $0736f
          29552 => x"80", -- $07370
          29553 => x"80", -- $07371
          29554 => x"80", -- $07372
          29555 => x"80", -- $07373
          29556 => x"80", -- $07374
          29557 => x"80", -- $07375
          29558 => x"80", -- $07376
          29559 => x"80", -- $07377
          29560 => x"7f", -- $07378
          29561 => x"7f", -- $07379
          29562 => x"7f", -- $0737a
          29563 => x"7f", -- $0737b
          29564 => x"7f", -- $0737c
          29565 => x"7f", -- $0737d
          29566 => x"7f", -- $0737e
          29567 => x"7f", -- $0737f
          29568 => x"7f", -- $07380
          29569 => x"7f", -- $07381
          29570 => x"7f", -- $07382
          29571 => x"7f", -- $07383
          29572 => x"7f", -- $07384
          29573 => x"7f", -- $07385
          29574 => x"7f", -- $07386
          29575 => x"7e", -- $07387
          29576 => x"7e", -- $07388
          29577 => x"7e", -- $07389
          29578 => x"7e", -- $0738a
          29579 => x"7e", -- $0738b
          29580 => x"7e", -- $0738c
          29581 => x"7e", -- $0738d
          29582 => x"7e", -- $0738e
          29583 => x"7f", -- $0738f
          29584 => x"7e", -- $07390
          29585 => x"7f", -- $07391
          29586 => x"7f", -- $07392
          29587 => x"7f", -- $07393
          29588 => x"7f", -- $07394
          29589 => x"7f", -- $07395
          29590 => x"7f", -- $07396
          29591 => x"7f", -- $07397
          29592 => x"7f", -- $07398
          29593 => x"7f", -- $07399
          29594 => x"7f", -- $0739a
          29595 => x"7f", -- $0739b
          29596 => x"7f", -- $0739c
          29597 => x"7f", -- $0739d
          29598 => x"7f", -- $0739e
          29599 => x"7e", -- $0739f
          29600 => x"7e", -- $073a0
          29601 => x"7e", -- $073a1
          29602 => x"7e", -- $073a2
          29603 => x"7e", -- $073a3
          29604 => x"7e", -- $073a4
          29605 => x"7e", -- $073a5
          29606 => x"7e", -- $073a6
          29607 => x"7e", -- $073a7
          29608 => x"7e", -- $073a8
          29609 => x"7e", -- $073a9
          29610 => x"7e", -- $073aa
          29611 => x"7e", -- $073ab
          29612 => x"7e", -- $073ac
          29613 => x"7e", -- $073ad
          29614 => x"7e", -- $073ae
          29615 => x"7e", -- $073af
          29616 => x"7e", -- $073b0
          29617 => x"7e", -- $073b1
          29618 => x"7e", -- $073b2
          29619 => x"7e", -- $073b3
          29620 => x"7e", -- $073b4
          29621 => x"7e", -- $073b5
          29622 => x"7e", -- $073b6
          29623 => x"7e", -- $073b7
          29624 => x"7d", -- $073b8
          29625 => x"7d", -- $073b9
          29626 => x"7d", -- $073ba
          29627 => x"7d", -- $073bb
          29628 => x"7d", -- $073bc
          29629 => x"7d", -- $073bd
          29630 => x"7e", -- $073be
          29631 => x"7d", -- $073bf
          29632 => x"7e", -- $073c0
          29633 => x"7e", -- $073c1
          29634 => x"7e", -- $073c2
          29635 => x"7e", -- $073c3
          29636 => x"7e", -- $073c4
          29637 => x"7e", -- $073c5
          29638 => x"7e", -- $073c6
          29639 => x"7e", -- $073c7
          29640 => x"7e", -- $073c8
          29641 => x"7e", -- $073c9
          29642 => x"7e", -- $073ca
          29643 => x"7e", -- $073cb
          29644 => x"7e", -- $073cc
          29645 => x"7e", -- $073cd
          29646 => x"7e", -- $073ce
          29647 => x"7e", -- $073cf
          29648 => x"7e", -- $073d0
          29649 => x"7e", -- $073d1
          29650 => x"7e", -- $073d2
          29651 => x"7e", -- $073d3
          29652 => x"7e", -- $073d4
          29653 => x"7e", -- $073d5
          29654 => x"7e", -- $073d6
          29655 => x"7e", -- $073d7
          29656 => x"7e", -- $073d8
          29657 => x"7e", -- $073d9
          29658 => x"7e", -- $073da
          29659 => x"7e", -- $073db
          29660 => x"7e", -- $073dc
          29661 => x"7e", -- $073dd
          29662 => x"7e", -- $073de
          29663 => x"7e", -- $073df
          29664 => x"7e", -- $073e0
          29665 => x"7e", -- $073e1
          29666 => x"7e", -- $073e2
          29667 => x"7e", -- $073e3
          29668 => x"7e", -- $073e4
          29669 => x"7e", -- $073e5
          29670 => x"7e", -- $073e6
          29671 => x"7e", -- $073e7
          29672 => x"7e", -- $073e8
          29673 => x"7d", -- $073e9
          29674 => x"7d", -- $073ea
          29675 => x"7d", -- $073eb
          29676 => x"7d", -- $073ec
          29677 => x"7d", -- $073ed
          29678 => x"7d", -- $073ee
          29679 => x"7d", -- $073ef
          29680 => x"7d", -- $073f0
          29681 => x"7d", -- $073f1
          29682 => x"7d", -- $073f2
          29683 => x"7e", -- $073f3
          29684 => x"7e", -- $073f4
          29685 => x"7e", -- $073f5
          29686 => x"7e", -- $073f6
          29687 => x"7e", -- $073f7
          29688 => x"7e", -- $073f8
          29689 => x"7e", -- $073f9
          29690 => x"7e", -- $073fa
          29691 => x"7e", -- $073fb
          29692 => x"7e", -- $073fc
          29693 => x"7e", -- $073fd
          29694 => x"7e", -- $073fe
          29695 => x"7e", -- $073ff
          29696 => x"7e", -- $07400
          29697 => x"7e", -- $07401
          29698 => x"7e", -- $07402
          29699 => x"7e", -- $07403
          29700 => x"7d", -- $07404
          29701 => x"7d", -- $07405
          29702 => x"7d", -- $07406
          29703 => x"7d", -- $07407
          29704 => x"7d", -- $07408
          29705 => x"7d", -- $07409
          29706 => x"7d", -- $0740a
          29707 => x"7d", -- $0740b
          29708 => x"7d", -- $0740c
          29709 => x"7d", -- $0740d
          29710 => x"7d", -- $0740e
          29711 => x"7d", -- $0740f
          29712 => x"7d", -- $07410
          29713 => x"7d", -- $07411
          29714 => x"7d", -- $07412
          29715 => x"7d", -- $07413
          29716 => x"7d", -- $07414
          29717 => x"7d", -- $07415
          29718 => x"7d", -- $07416
          29719 => x"7d", -- $07417
          29720 => x"7d", -- $07418
          29721 => x"7d", -- $07419
          29722 => x"7d", -- $0741a
          29723 => x"7d", -- $0741b
          29724 => x"7d", -- $0741c
          29725 => x"7d", -- $0741d
          29726 => x"7d", -- $0741e
          29727 => x"7d", -- $0741f
          29728 => x"7d", -- $07420
          29729 => x"7d", -- $07421
          29730 => x"7d", -- $07422
          29731 => x"7d", -- $07423
          29732 => x"7d", -- $07424
          29733 => x"7d", -- $07425
          29734 => x"7d", -- $07426
          29735 => x"7d", -- $07427
          29736 => x"7d", -- $07428
          29737 => x"7d", -- $07429
          29738 => x"7d", -- $0742a
          29739 => x"7d", -- $0742b
          29740 => x"7d", -- $0742c
          29741 => x"7d", -- $0742d
          29742 => x"7d", -- $0742e
          29743 => x"7d", -- $0742f
          29744 => x"7d", -- $07430
          29745 => x"7d", -- $07431
          29746 => x"7d", -- $07432
          29747 => x"7d", -- $07433
          29748 => x"7d", -- $07434
          29749 => x"7d", -- $07435
          29750 => x"7d", -- $07436
          29751 => x"7d", -- $07437
          29752 => x"7d", -- $07438
          29753 => x"7d", -- $07439
          29754 => x"7d", -- $0743a
          29755 => x"7d", -- $0743b
          29756 => x"7d", -- $0743c
          29757 => x"7d", -- $0743d
          29758 => x"7d", -- $0743e
          29759 => x"7d", -- $0743f
          29760 => x"7d", -- $07440
          29761 => x"7d", -- $07441
          29762 => x"7d", -- $07442
          29763 => x"7d", -- $07443
          29764 => x"7d", -- $07444
          29765 => x"7d", -- $07445
          29766 => x"7d", -- $07446
          29767 => x"7d", -- $07447
          29768 => x"7d", -- $07448
          29769 => x"7d", -- $07449
          29770 => x"7d", -- $0744a
          29771 => x"7d", -- $0744b
          29772 => x"7d", -- $0744c
          29773 => x"7d", -- $0744d
          29774 => x"7e", -- $0744e
          29775 => x"7e", -- $0744f
          29776 => x"7e", -- $07450
          29777 => x"7e", -- $07451
          29778 => x"7e", -- $07452
          29779 => x"7e", -- $07453
          29780 => x"7e", -- $07454
          29781 => x"7e", -- $07455
          29782 => x"7e", -- $07456
          29783 => x"7e", -- $07457
          29784 => x"7e", -- $07458
          29785 => x"7e", -- $07459
          29786 => x"7e", -- $0745a
          29787 => x"7e", -- $0745b
          29788 => x"7e", -- $0745c
          29789 => x"7e", -- $0745d
          29790 => x"7e", -- $0745e
          29791 => x"7e", -- $0745f
          29792 => x"7e", -- $07460
          29793 => x"7e", -- $07461
          29794 => x"7e", -- $07462
          29795 => x"7e", -- $07463
          29796 => x"7e", -- $07464
          29797 => x"7e", -- $07465
          29798 => x"7e", -- $07466
          29799 => x"7e", -- $07467
          29800 => x"7e", -- $07468
          29801 => x"7e", -- $07469
          29802 => x"7e", -- $0746a
          29803 => x"7e", -- $0746b
          29804 => x"7e", -- $0746c
          29805 => x"7e", -- $0746d
          29806 => x"7e", -- $0746e
          29807 => x"7e", -- $0746f
          29808 => x"7e", -- $07470
          29809 => x"7e", -- $07471
          29810 => x"7e", -- $07472
          29811 => x"7e", -- $07473
          29812 => x"7e", -- $07474
          29813 => x"7e", -- $07475
          29814 => x"7e", -- $07476
          29815 => x"7e", -- $07477
          29816 => x"7e", -- $07478
          29817 => x"7f", -- $07479
          29818 => x"7f", -- $0747a
          29819 => x"7f", -- $0747b
          29820 => x"7f", -- $0747c
          29821 => x"7f", -- $0747d
          29822 => x"7f", -- $0747e
          29823 => x"7f", -- $0747f
          29824 => x"7f", -- $07480
          29825 => x"7f", -- $07481
          29826 => x"7f", -- $07482
          29827 => x"7e", -- $07483
          29828 => x"7e", -- $07484
          29829 => x"7e", -- $07485
          29830 => x"7e", -- $07486
          29831 => x"7e", -- $07487
          29832 => x"7e", -- $07488
          29833 => x"7e", -- $07489
          29834 => x"7e", -- $0748a
          29835 => x"7e", -- $0748b
          29836 => x"7e", -- $0748c
          29837 => x"7e", -- $0748d
          29838 => x"7e", -- $0748e
          29839 => x"7e", -- $0748f
          29840 => x"7e", -- $07490
          29841 => x"7e", -- $07491
          29842 => x"7e", -- $07492
          29843 => x"7e", -- $07493
          29844 => x"7e", -- $07494
          29845 => x"7e", -- $07495
          29846 => x"7e", -- $07496
          29847 => x"7e", -- $07497
          29848 => x"7e", -- $07498
          29849 => x"7e", -- $07499
          29850 => x"7e", -- $0749a
          29851 => x"7e", -- $0749b
          29852 => x"7f", -- $0749c
          29853 => x"7f", -- $0749d
          29854 => x"7f", -- $0749e
          29855 => x"7f", -- $0749f
          29856 => x"7f", -- $074a0
          29857 => x"7f", -- $074a1
          29858 => x"7f", -- $074a2
          29859 => x"7f", -- $074a3
          29860 => x"7f", -- $074a4
          29861 => x"7f", -- $074a5
          29862 => x"7f", -- $074a6
          29863 => x"7f", -- $074a7
          29864 => x"7f", -- $074a8
          29865 => x"7f", -- $074a9
          29866 => x"7f", -- $074aa
          29867 => x"7f", -- $074ab
          29868 => x"7f", -- $074ac
          29869 => x"7f", -- $074ad
          29870 => x"7f", -- $074ae
          29871 => x"7f", -- $074af
          29872 => x"7f", -- $074b0
          29873 => x"7f", -- $074b1
          29874 => x"7f", -- $074b2
          29875 => x"7f", -- $074b3
          29876 => x"7f", -- $074b4
          29877 => x"7f", -- $074b5
          29878 => x"7f", -- $074b6
          29879 => x"7f", -- $074b7
          29880 => x"7f", -- $074b8
          29881 => x"7f", -- $074b9
          29882 => x"7f", -- $074ba
          29883 => x"7f", -- $074bb
          29884 => x"7f", -- $074bc
          29885 => x"7f", -- $074bd
          29886 => x"7f", -- $074be
          29887 => x"7f", -- $074bf
          29888 => x"7f", -- $074c0
          29889 => x"7f", -- $074c1
          29890 => x"7f", -- $074c2
          29891 => x"7f", -- $074c3
          29892 => x"80", -- $074c4
          29893 => x"80", -- $074c5
          29894 => x"80", -- $074c6
          29895 => x"80", -- $074c7
          29896 => x"80", -- $074c8
          29897 => x"80", -- $074c9
          29898 => x"80", -- $074ca
          29899 => x"80", -- $074cb
          29900 => x"80", -- $074cc
          29901 => x"80", -- $074cd
          29902 => x"80", -- $074ce
          29903 => x"80", -- $074cf
          29904 => x"80", -- $074d0
          29905 => x"80", -- $074d1
          29906 => x"80", -- $074d2
          29907 => x"80", -- $074d3
          29908 => x"80", -- $074d4
          29909 => x"80", -- $074d5
          29910 => x"80", -- $074d6
          29911 => x"80", -- $074d7
          29912 => x"80", -- $074d8
          29913 => x"80", -- $074d9
          29914 => x"80", -- $074da
          29915 => x"80", -- $074db
          29916 => x"80", -- $074dc
          29917 => x"80", -- $074dd
          29918 => x"80", -- $074de
          29919 => x"80", -- $074df
          29920 => x"80", -- $074e0
          29921 => x"80", -- $074e1
          29922 => x"80", -- $074e2
          29923 => x"80", -- $074e3
          29924 => x"80", -- $074e4
          29925 => x"80", -- $074e5
          29926 => x"80", -- $074e6
          29927 => x"80", -- $074e7
          29928 => x"80", -- $074e8
          29929 => x"80", -- $074e9
          29930 => x"80", -- $074ea
          29931 => x"80", -- $074eb
          29932 => x"80", -- $074ec
          29933 => x"80", -- $074ed
          29934 => x"80", -- $074ee
          29935 => x"80", -- $074ef
          29936 => x"80", -- $074f0
          29937 => x"80", -- $074f1
          29938 => x"80", -- $074f2
          29939 => x"80", -- $074f3
          29940 => x"80", -- $074f4
          29941 => x"80", -- $074f5
          29942 => x"80", -- $074f6
          29943 => x"80", -- $074f7
          29944 => x"80", -- $074f8
          29945 => x"80", -- $074f9
          29946 => x"80", -- $074fa
          29947 => x"80", -- $074fb
          29948 => x"80", -- $074fc
          29949 => x"80", -- $074fd
          29950 => x"80", -- $074fe
          29951 => x"80", -- $074ff
          29952 => x"80", -- $07500
          29953 => x"80", -- $07501
          29954 => x"80", -- $07502
          29955 => x"80", -- $07503
          29956 => x"80", -- $07504
          29957 => x"80", -- $07505
          29958 => x"80", -- $07506
          29959 => x"80", -- $07507
          29960 => x"80", -- $07508
          29961 => x"80", -- $07509
          29962 => x"80", -- $0750a
          29963 => x"80", -- $0750b
          29964 => x"80", -- $0750c
          29965 => x"80", -- $0750d
          29966 => x"80", -- $0750e
          29967 => x"80", -- $0750f
          29968 => x"80", -- $07510
          29969 => x"80", -- $07511
          29970 => x"80", -- $07512
          29971 => x"80", -- $07513
          29972 => x"81", -- $07514
          29973 => x"81", -- $07515
          29974 => x"81", -- $07516
          29975 => x"81", -- $07517
          29976 => x"81", -- $07518
          29977 => x"81", -- $07519
          29978 => x"81", -- $0751a
          29979 => x"81", -- $0751b
          29980 => x"81", -- $0751c
          29981 => x"81", -- $0751d
          29982 => x"81", -- $0751e
          29983 => x"81", -- $0751f
          29984 => x"81", -- $07520
          29985 => x"81", -- $07521
          29986 => x"81", -- $07522
          29987 => x"81", -- $07523
          29988 => x"81", -- $07524
          29989 => x"81", -- $07525
          29990 => x"81", -- $07526
          29991 => x"81", -- $07527
          29992 => x"81", -- $07528
          29993 => x"81", -- $07529
          29994 => x"81", -- $0752a
          29995 => x"81", -- $0752b
          29996 => x"81", -- $0752c
          29997 => x"81", -- $0752d
          29998 => x"81", -- $0752e
          29999 => x"81", -- $0752f
          30000 => x"81", -- $07530
          30001 => x"81", -- $07531
          30002 => x"81", -- $07532
          30003 => x"81", -- $07533
          30004 => x"81", -- $07534
          30005 => x"81", -- $07535
          30006 => x"81", -- $07536
          30007 => x"81", -- $07537
          30008 => x"81", -- $07538
          30009 => x"81", -- $07539
          30010 => x"81", -- $0753a
          30011 => x"81", -- $0753b
          30012 => x"81", -- $0753c
          30013 => x"81", -- $0753d
          30014 => x"82", -- $0753e
          30015 => x"82", -- $0753f
          30016 => x"82", -- $07540
          30017 => x"82", -- $07541
          30018 => x"82", -- $07542
          30019 => x"82", -- $07543
          30020 => x"82", -- $07544
          30021 => x"82", -- $07545
          30022 => x"82", -- $07546
          30023 => x"82", -- $07547
          30024 => x"82", -- $07548
          30025 => x"81", -- $07549
          30026 => x"81", -- $0754a
          30027 => x"81", -- $0754b
          30028 => x"81", -- $0754c
          30029 => x"82", -- $0754d
          30030 => x"82", -- $0754e
          30031 => x"82", -- $0754f
          30032 => x"82", -- $07550
          30033 => x"82", -- $07551
          30034 => x"82", -- $07552
          30035 => x"82", -- $07553
          30036 => x"82", -- $07554
          30037 => x"82", -- $07555
          30038 => x"82", -- $07556
          30039 => x"82", -- $07557
          30040 => x"82", -- $07558
          30041 => x"82", -- $07559
          30042 => x"82", -- $0755a
          30043 => x"82", -- $0755b
          30044 => x"82", -- $0755c
          30045 => x"82", -- $0755d
          30046 => x"82", -- $0755e
          30047 => x"82", -- $0755f
          30048 => x"82", -- $07560
          30049 => x"83", -- $07561
          30050 => x"83", -- $07562
          30051 => x"83", -- $07563
          30052 => x"83", -- $07564
          30053 => x"83", -- $07565
          30054 => x"83", -- $07566
          30055 => x"83", -- $07567
          30056 => x"83", -- $07568
          30057 => x"83", -- $07569
          30058 => x"83", -- $0756a
          30059 => x"83", -- $0756b
          30060 => x"83", -- $0756c
          30061 => x"83", -- $0756d
          30062 => x"83", -- $0756e
          30063 => x"83", -- $0756f
          30064 => x"83", -- $07570
          30065 => x"83", -- $07571
          30066 => x"82", -- $07572
          30067 => x"82", -- $07573
          30068 => x"83", -- $07574
          30069 => x"83", -- $07575
          30070 => x"83", -- $07576
          30071 => x"83", -- $07577
          30072 => x"83", -- $07578
          30073 => x"83", -- $07579
          30074 => x"84", -- $0757a
          30075 => x"84", -- $0757b
          30076 => x"84", -- $0757c
          30077 => x"84", -- $0757d
          30078 => x"84", -- $0757e
          30079 => x"84", -- $0757f
          30080 => x"84", -- $07580
          30081 => x"84", -- $07581
          30082 => x"84", -- $07582
          30083 => x"84", -- $07583
          30084 => x"84", -- $07584
          30085 => x"84", -- $07585
          30086 => x"84", -- $07586
          30087 => x"84", -- $07587
          30088 => x"84", -- $07588
          30089 => x"84", -- $07589
          30090 => x"84", -- $0758a
          30091 => x"84", -- $0758b
          30092 => x"84", -- $0758c
          30093 => x"84", -- $0758d
          30094 => x"84", -- $0758e
          30095 => x"84", -- $0758f
          30096 => x"84", -- $07590
          30097 => x"84", -- $07591
          30098 => x"84", -- $07592
          30099 => x"84", -- $07593
          30100 => x"84", -- $07594
          30101 => x"83", -- $07595
          30102 => x"83", -- $07596
          30103 => x"84", -- $07597
          30104 => x"84", -- $07598
          30105 => x"83", -- $07599
          30106 => x"83", -- $0759a
          30107 => x"83", -- $0759b
          30108 => x"84", -- $0759c
          30109 => x"84", -- $0759d
          30110 => x"84", -- $0759e
          30111 => x"84", -- $0759f
          30112 => x"84", -- $075a0
          30113 => x"84", -- $075a1
          30114 => x"84", -- $075a2
          30115 => x"84", -- $075a3
          30116 => x"85", -- $075a4
          30117 => x"85", -- $075a5
          30118 => x"85", -- $075a6
          30119 => x"85", -- $075a7
          30120 => x"85", -- $075a8
          30121 => x"85", -- $075a9
          30122 => x"84", -- $075aa
          30123 => x"84", -- $075ab
          30124 => x"84", -- $075ac
          30125 => x"84", -- $075ad
          30126 => x"84", -- $075ae
          30127 => x"84", -- $075af
          30128 => x"84", -- $075b0
          30129 => x"84", -- $075b1
          30130 => x"83", -- $075b2
          30131 => x"83", -- $075b3
          30132 => x"83", -- $075b4
          30133 => x"83", -- $075b5
          30134 => x"83", -- $075b6
          30135 => x"83", -- $075b7
          30136 => x"83", -- $075b8
          30137 => x"83", -- $075b9
          30138 => x"83", -- $075ba
          30139 => x"83", -- $075bb
          30140 => x"83", -- $075bc
          30141 => x"83", -- $075bd
          30142 => x"83", -- $075be
          30143 => x"83", -- $075bf
          30144 => x"83", -- $075c0
          30145 => x"83", -- $075c1
          30146 => x"83", -- $075c2
          30147 => x"83", -- $075c3
          30148 => x"83", -- $075c4
          30149 => x"83", -- $075c5
          30150 => x"83", -- $075c6
          30151 => x"83", -- $075c7
          30152 => x"83", -- $075c8
          30153 => x"83", -- $075c9
          30154 => x"83", -- $075ca
          30155 => x"83", -- $075cb
          30156 => x"83", -- $075cc
          30157 => x"83", -- $075cd
          30158 => x"83", -- $075ce
          30159 => x"83", -- $075cf
          30160 => x"83", -- $075d0
          30161 => x"83", -- $075d1
          30162 => x"83", -- $075d2
          30163 => x"82", -- $075d3
          30164 => x"82", -- $075d4
          30165 => x"82", -- $075d5
          30166 => x"82", -- $075d6
          30167 => x"82", -- $075d7
          30168 => x"82", -- $075d8
          30169 => x"81", -- $075d9
          30170 => x"81", -- $075da
          30171 => x"81", -- $075db
          30172 => x"81", -- $075dc
          30173 => x"81", -- $075dd
          30174 => x"81", -- $075de
          30175 => x"81", -- $075df
          30176 => x"81", -- $075e0
          30177 => x"81", -- $075e1
          30178 => x"81", -- $075e2
          30179 => x"81", -- $075e3
          30180 => x"81", -- $075e4
          30181 => x"81", -- $075e5
          30182 => x"81", -- $075e6
          30183 => x"81", -- $075e7
          30184 => x"82", -- $075e8
          30185 => x"82", -- $075e9
          30186 => x"82", -- $075ea
          30187 => x"82", -- $075eb
          30188 => x"82", -- $075ec
          30189 => x"82", -- $075ed
          30190 => x"82", -- $075ee
          30191 => x"82", -- $075ef
          30192 => x"82", -- $075f0
          30193 => x"82", -- $075f1
          30194 => x"82", -- $075f2
          30195 => x"82", -- $075f3
          30196 => x"82", -- $075f4
          30197 => x"82", -- $075f5
          30198 => x"81", -- $075f6
          30199 => x"81", -- $075f7
          30200 => x"81", -- $075f8
          30201 => x"81", -- $075f9
          30202 => x"81", -- $075fa
          30203 => x"81", -- $075fb
          30204 => x"81", -- $075fc
          30205 => x"80", -- $075fd
          30206 => x"81", -- $075fe
          30207 => x"80", -- $075ff
          30208 => x"80", -- $07600
          30209 => x"80", -- $07601
          30210 => x"80", -- $07602
          30211 => x"80", -- $07603
          30212 => x"80", -- $07604
          30213 => x"80", -- $07605
          30214 => x"80", -- $07606
          30215 => x"80", -- $07607
          30216 => x"80", -- $07608
          30217 => x"81", -- $07609
          30218 => x"81", -- $0760a
          30219 => x"81", -- $0760b
          30220 => x"81", -- $0760c
          30221 => x"81", -- $0760d
          30222 => x"81", -- $0760e
          30223 => x"81", -- $0760f
          30224 => x"82", -- $07610
          30225 => x"82", -- $07611
          30226 => x"82", -- $07612
          30227 => x"82", -- $07613
          30228 => x"82", -- $07614
          30229 => x"82", -- $07615
          30230 => x"82", -- $07616
          30231 => x"82", -- $07617
          30232 => x"81", -- $07618
          30233 => x"81", -- $07619
          30234 => x"81", -- $0761a
          30235 => x"81", -- $0761b
          30236 => x"81", -- $0761c
          30237 => x"81", -- $0761d
          30238 => x"81", -- $0761e
          30239 => x"80", -- $0761f
          30240 => x"80", -- $07620
          30241 => x"80", -- $07621
          30242 => x"80", -- $07622
          30243 => x"80", -- $07623
          30244 => x"80", -- $07624
          30245 => x"80", -- $07625
          30246 => x"80", -- $07626
          30247 => x"80", -- $07627
          30248 => x"80", -- $07628
          30249 => x"80", -- $07629
          30250 => x"80", -- $0762a
          30251 => x"80", -- $0762b
          30252 => x"80", -- $0762c
          30253 => x"80", -- $0762d
          30254 => x"80", -- $0762e
          30255 => x"81", -- $0762f
          30256 => x"81", -- $07630
          30257 => x"81", -- $07631
          30258 => x"81", -- $07632
          30259 => x"81", -- $07633
          30260 => x"81", -- $07634
          30261 => x"81", -- $07635
          30262 => x"82", -- $07636
          30263 => x"82", -- $07637
          30264 => x"82", -- $07638
          30265 => x"81", -- $07639
          30266 => x"82", -- $0763a
          30267 => x"82", -- $0763b
          30268 => x"81", -- $0763c
          30269 => x"81", -- $0763d
          30270 => x"81", -- $0763e
          30271 => x"81", -- $0763f
          30272 => x"80", -- $07640
          30273 => x"80", -- $07641
          30274 => x"80", -- $07642
          30275 => x"80", -- $07643
          30276 => x"80", -- $07644
          30277 => x"80", -- $07645
          30278 => x"80", -- $07646
          30279 => x"80", -- $07647
          30280 => x"80", -- $07648
          30281 => x"80", -- $07649
          30282 => x"80", -- $0764a
          30283 => x"80", -- $0764b
          30284 => x"80", -- $0764c
          30285 => x"80", -- $0764d
          30286 => x"80", -- $0764e
          30287 => x"80", -- $0764f
          30288 => x"80", -- $07650
          30289 => x"80", -- $07651
          30290 => x"80", -- $07652
          30291 => x"80", -- $07653
          30292 => x"80", -- $07654
          30293 => x"80", -- $07655
          30294 => x"81", -- $07656
          30295 => x"81", -- $07657
          30296 => x"81", -- $07658
          30297 => x"81", -- $07659
          30298 => x"81", -- $0765a
          30299 => x"81", -- $0765b
          30300 => x"81", -- $0765c
          30301 => x"81", -- $0765d
          30302 => x"81", -- $0765e
          30303 => x"81", -- $0765f
          30304 => x"81", -- $07660
          30305 => x"80", -- $07661
          30306 => x"80", -- $07662
          30307 => x"80", -- $07663
          30308 => x"80", -- $07664
          30309 => x"80", -- $07665
          30310 => x"80", -- $07666
          30311 => x"80", -- $07667
          30312 => x"80", -- $07668
          30313 => x"80", -- $07669
          30314 => x"7f", -- $0766a
          30315 => x"80", -- $0766b
          30316 => x"7f", -- $0766c
          30317 => x"7f", -- $0766d
          30318 => x"7f", -- $0766e
          30319 => x"7f", -- $0766f
          30320 => x"7f", -- $07670
          30321 => x"7f", -- $07671
          30322 => x"80", -- $07672
          30323 => x"80", -- $07673
          30324 => x"80", -- $07674
          30325 => x"80", -- $07675
          30326 => x"80", -- $07676
          30327 => x"80", -- $07677
          30328 => x"80", -- $07678
          30329 => x"80", -- $07679
          30330 => x"80", -- $0767a
          30331 => x"80", -- $0767b
          30332 => x"80", -- $0767c
          30333 => x"80", -- $0767d
          30334 => x"80", -- $0767e
          30335 => x"80", -- $0767f
          30336 => x"80", -- $07680
          30337 => x"80", -- $07681
          30338 => x"80", -- $07682
          30339 => x"80", -- $07683
          30340 => x"80", -- $07684
          30341 => x"80", -- $07685
          30342 => x"80", -- $07686
          30343 => x"80", -- $07687
          30344 => x"80", -- $07688
          30345 => x"7f", -- $07689
          30346 => x"7f", -- $0768a
          30347 => x"7f", -- $0768b
          30348 => x"7f", -- $0768c
          30349 => x"7f", -- $0768d
          30350 => x"7f", -- $0768e
          30351 => x"7f", -- $0768f
          30352 => x"7f", -- $07690
          30353 => x"7e", -- $07691
          30354 => x"7e", -- $07692
          30355 => x"7e", -- $07693
          30356 => x"7e", -- $07694
          30357 => x"7e", -- $07695
          30358 => x"7f", -- $07696
          30359 => x"7f", -- $07697
          30360 => x"7f", -- $07698
          30361 => x"7f", -- $07699
          30362 => x"7f", -- $0769a
          30363 => x"7f", -- $0769b
          30364 => x"7f", -- $0769c
          30365 => x"80", -- $0769d
          30366 => x"80", -- $0769e
          30367 => x"7f", -- $0769f
          30368 => x"80", -- $076a0
          30369 => x"80", -- $076a1
          30370 => x"80", -- $076a2
          30371 => x"80", -- $076a3
          30372 => x"80", -- $076a4
          30373 => x"80", -- $076a5
          30374 => x"80", -- $076a6
          30375 => x"80", -- $076a7
          30376 => x"80", -- $076a8
          30377 => x"7f", -- $076a9
          30378 => x"7f", -- $076aa
          30379 => x"7f", -- $076ab
          30380 => x"7f", -- $076ac
          30381 => x"7e", -- $076ad
          30382 => x"7e", -- $076ae
          30383 => x"7e", -- $076af
          30384 => x"7e", -- $076b0
          30385 => x"7e", -- $076b1
          30386 => x"7e", -- $076b2
          30387 => x"7e", -- $076b3
          30388 => x"7e", -- $076b4
          30389 => x"7e", -- $076b5
          30390 => x"7e", -- $076b6
          30391 => x"7e", -- $076b7
          30392 => x"7e", -- $076b8
          30393 => x"7e", -- $076b9
          30394 => x"7e", -- $076ba
          30395 => x"7e", -- $076bb
          30396 => x"7e", -- $076bc
          30397 => x"7e", -- $076bd
          30398 => x"7e", -- $076be
          30399 => x"7e", -- $076bf
          30400 => x"7e", -- $076c0
          30401 => x"7f", -- $076c1
          30402 => x"7f", -- $076c2
          30403 => x"7f", -- $076c3
          30404 => x"7f", -- $076c4
          30405 => x"7f", -- $076c5
          30406 => x"7f", -- $076c6
          30407 => x"7f", -- $076c7
          30408 => x"7f", -- $076c8
          30409 => x"7f", -- $076c9
          30410 => x"7f", -- $076ca
          30411 => x"7f", -- $076cb
          30412 => x"7f", -- $076cc
          30413 => x"7e", -- $076cd
          30414 => x"7e", -- $076ce
          30415 => x"7e", -- $076cf
          30416 => x"7e", -- $076d0
          30417 => x"7e", -- $076d1
          30418 => x"7e", -- $076d2
          30419 => x"7d", -- $076d3
          30420 => x"7d", -- $076d4
          30421 => x"7d", -- $076d5
          30422 => x"7d", -- $076d6
          30423 => x"7d", -- $076d7
          30424 => x"7c", -- $076d8
          30425 => x"7d", -- $076d9
          30426 => x"7d", -- $076da
          30427 => x"7d", -- $076db
          30428 => x"7d", -- $076dc
          30429 => x"7d", -- $076dd
          30430 => x"7d", -- $076de
          30431 => x"7d", -- $076df
          30432 => x"7d", -- $076e0
          30433 => x"7e", -- $076e1
          30434 => x"7e", -- $076e2
          30435 => x"7e", -- $076e3
          30436 => x"7e", -- $076e4
          30437 => x"7e", -- $076e5
          30438 => x"7e", -- $076e6
          30439 => x"7e", -- $076e7
          30440 => x"7f", -- $076e8
          30441 => x"7f", -- $076e9
          30442 => x"7e", -- $076ea
          30443 => x"7f", -- $076eb
          30444 => x"7f", -- $076ec
          30445 => x"7e", -- $076ed
          30446 => x"7e", -- $076ee
          30447 => x"7e", -- $076ef
          30448 => x"7e", -- $076f0
          30449 => x"7d", -- $076f1
          30450 => x"7d", -- $076f2
          30451 => x"7d", -- $076f3
          30452 => x"7d", -- $076f4
          30453 => x"7d", -- $076f5
          30454 => x"7d", -- $076f6
          30455 => x"7d", -- $076f7
          30456 => x"7c", -- $076f8
          30457 => x"7c", -- $076f9
          30458 => x"7c", -- $076fa
          30459 => x"7c", -- $076fb
          30460 => x"7c", -- $076fc
          30461 => x"7c", -- $076fd
          30462 => x"7c", -- $076fe
          30463 => x"7c", -- $076ff
          30464 => x"7d", -- $07700
          30465 => x"7d", -- $07701
          30466 => x"7d", -- $07702
          30467 => x"7d", -- $07703
          30468 => x"7d", -- $07704
          30469 => x"7d", -- $07705
          30470 => x"7d", -- $07706
          30471 => x"7e", -- $07707
          30472 => x"7e", -- $07708
          30473 => x"7e", -- $07709
          30474 => x"7e", -- $0770a
          30475 => x"7e", -- $0770b
          30476 => x"7e", -- $0770c
          30477 => x"7e", -- $0770d
          30478 => x"7e", -- $0770e
          30479 => x"7f", -- $0770f
          30480 => x"7f", -- $07710
          30481 => x"7f", -- $07711
          30482 => x"7e", -- $07712
          30483 => x"7e", -- $07713
          30484 => x"7e", -- $07714
          30485 => x"7e", -- $07715
          30486 => x"7e", -- $07716
          30487 => x"7e", -- $07717
          30488 => x"7d", -- $07718
          30489 => x"7d", -- $07719
          30490 => x"7d", -- $0771a
          30491 => x"7d", -- $0771b
          30492 => x"7d", -- $0771c
          30493 => x"7d", -- $0771d
          30494 => x"7d", -- $0771e
          30495 => x"7d", -- $0771f
          30496 => x"7d", -- $07720
          30497 => x"7d", -- $07721
          30498 => x"7d", -- $07722
          30499 => x"7d", -- $07723
          30500 => x"7d", -- $07724
          30501 => x"7d", -- $07725
          30502 => x"7d", -- $07726
          30503 => x"7d", -- $07727
          30504 => x"7e", -- $07728
          30505 => x"7e", -- $07729
          30506 => x"7e", -- $0772a
          30507 => x"7e", -- $0772b
          30508 => x"7e", -- $0772c
          30509 => x"7e", -- $0772d
          30510 => x"7e", -- $0772e
          30511 => x"7e", -- $0772f
          30512 => x"7f", -- $07730
          30513 => x"7f", -- $07731
          30514 => x"7f", -- $07732
          30515 => x"7f", -- $07733
          30516 => x"7f", -- $07734
          30517 => x"7f", -- $07735
          30518 => x"7f", -- $07736
          30519 => x"7e", -- $07737
          30520 => x"7e", -- $07738
          30521 => x"7e", -- $07739
          30522 => x"7e", -- $0773a
          30523 => x"7e", -- $0773b
          30524 => x"7d", -- $0773c
          30525 => x"7d", -- $0773d
          30526 => x"7d", -- $0773e
          30527 => x"7d", -- $0773f
          30528 => x"7d", -- $07740
          30529 => x"7d", -- $07741
          30530 => x"7d", -- $07742
          30531 => x"7d", -- $07743
          30532 => x"7d", -- $07744
          30533 => x"7d", -- $07745
          30534 => x"7d", -- $07746
          30535 => x"7d", -- $07747
          30536 => x"7d", -- $07748
          30537 => x"7e", -- $07749
          30538 => x"7e", -- $0774a
          30539 => x"7e", -- $0774b
          30540 => x"7e", -- $0774c
          30541 => x"7e", -- $0774d
          30542 => x"7e", -- $0774e
          30543 => x"7e", -- $0774f
          30544 => x"7f", -- $07750
          30545 => x"7f", -- $07751
          30546 => x"7f", -- $07752
          30547 => x"7f", -- $07753
          30548 => x"7f", -- $07754
          30549 => x"7f", -- $07755
          30550 => x"7f", -- $07756
          30551 => x"80", -- $07757
          30552 => x"7f", -- $07758
          30553 => x"7f", -- $07759
          30554 => x"7f", -- $0775a
          30555 => x"7f", -- $0775b
          30556 => x"7f", -- $0775c
          30557 => x"7f", -- $0775d
          30558 => x"7e", -- $0775e
          30559 => x"7e", -- $0775f
          30560 => x"7e", -- $07760
          30561 => x"7e", -- $07761
          30562 => x"7e", -- $07762
          30563 => x"7e", -- $07763
          30564 => x"7e", -- $07764
          30565 => x"7e", -- $07765
          30566 => x"7e", -- $07766
          30567 => x"7e", -- $07767
          30568 => x"7e", -- $07768
          30569 => x"7e", -- $07769
          30570 => x"7e", -- $0776a
          30571 => x"7e", -- $0776b
          30572 => x"7e", -- $0776c
          30573 => x"7e", -- $0776d
          30574 => x"7e", -- $0776e
          30575 => x"7e", -- $0776f
          30576 => x"7f", -- $07770
          30577 => x"7f", -- $07771
          30578 => x"7f", -- $07772
          30579 => x"7f", -- $07773
          30580 => x"7f", -- $07774
          30581 => x"7f", -- $07775
          30582 => x"7f", -- $07776
          30583 => x"7f", -- $07777
          30584 => x"80", -- $07778
          30585 => x"80", -- $07779
          30586 => x"80", -- $0777a
          30587 => x"80", -- $0777b
          30588 => x"80", -- $0777c
          30589 => x"80", -- $0777d
          30590 => x"7f", -- $0777e
          30591 => x"7f", -- $0777f
          30592 => x"7f", -- $07780
          30593 => x"7f", -- $07781
          30594 => x"7f", -- $07782
          30595 => x"7f", -- $07783
          30596 => x"7e", -- $07784
          30597 => x"7e", -- $07785
          30598 => x"7e", -- $07786
          30599 => x"7e", -- $07787
          30600 => x"7e", -- $07788
          30601 => x"7e", -- $07789
          30602 => x"7e", -- $0778a
          30603 => x"7e", -- $0778b
          30604 => x"7e", -- $0778c
          30605 => x"7e", -- $0778d
          30606 => x"7e", -- $0778e
          30607 => x"7e", -- $0778f
          30608 => x"7e", -- $07790
          30609 => x"7e", -- $07791
          30610 => x"7e", -- $07792
          30611 => x"7e", -- $07793
          30612 => x"7e", -- $07794
          30613 => x"7f", -- $07795
          30614 => x"7f", -- $07796
          30615 => x"7f", -- $07797
          30616 => x"7f", -- $07798
          30617 => x"7f", -- $07799
          30618 => x"7f", -- $0779a
          30619 => x"7f", -- $0779b
          30620 => x"7f", -- $0779c
          30621 => x"80", -- $0779d
          30622 => x"80", -- $0779e
          30623 => x"80", -- $0779f
          30624 => x"80", -- $077a0
          30625 => x"7f", -- $077a1
          30626 => x"7f", -- $077a2
          30627 => x"7f", -- $077a3
          30628 => x"7f", -- $077a4
          30629 => x"7f", -- $077a5
          30630 => x"7f", -- $077a6
          30631 => x"7e", -- $077a7
          30632 => x"7e", -- $077a8
          30633 => x"7e", -- $077a9
          30634 => x"7e", -- $077aa
          30635 => x"7e", -- $077ab
          30636 => x"7e", -- $077ac
          30637 => x"7e", -- $077ad
          30638 => x"7e", -- $077ae
          30639 => x"7e", -- $077af
          30640 => x"7e", -- $077b0
          30641 => x"7e", -- $077b1
          30642 => x"7e", -- $077b2
          30643 => x"7e", -- $077b3
          30644 => x"7e", -- $077b4
          30645 => x"7e", -- $077b5
          30646 => x"7e", -- $077b6
          30647 => x"7f", -- $077b7
          30648 => x"7f", -- $077b8
          30649 => x"7f", -- $077b9
          30650 => x"7f", -- $077ba
          30651 => x"7f", -- $077bb
          30652 => x"80", -- $077bc
          30653 => x"80", -- $077bd
          30654 => x"80", -- $077be
          30655 => x"80", -- $077bf
          30656 => x"80", -- $077c0
          30657 => x"80", -- $077c1
          30658 => x"80", -- $077c2
          30659 => x"80", -- $077c3
          30660 => x"80", -- $077c4
          30661 => x"80", -- $077c5
          30662 => x"80", -- $077c6
          30663 => x"80", -- $077c7
          30664 => x"80", -- $077c8
          30665 => x"80", -- $077c9
          30666 => x"80", -- $077ca
          30667 => x"7f", -- $077cb
          30668 => x"7f", -- $077cc
          30669 => x"7f", -- $077cd
          30670 => x"7f", -- $077ce
          30671 => x"7f", -- $077cf
          30672 => x"7f", -- $077d0
          30673 => x"7f", -- $077d1
          30674 => x"7f", -- $077d2
          30675 => x"7f", -- $077d3
          30676 => x"7f", -- $077d4
          30677 => x"7f", -- $077d5
          30678 => x"7f", -- $077d6
          30679 => x"7f", -- $077d7
          30680 => x"7f", -- $077d8
          30681 => x"7f", -- $077d9
          30682 => x"80", -- $077da
          30683 => x"80", -- $077db
          30684 => x"80", -- $077dc
          30685 => x"80", -- $077dd
          30686 => x"80", -- $077de
          30687 => x"80", -- $077df
          30688 => x"80", -- $077e0
          30689 => x"80", -- $077e1
          30690 => x"80", -- $077e2
          30691 => x"80", -- $077e3
          30692 => x"80", -- $077e4
          30693 => x"81", -- $077e5
          30694 => x"81", -- $077e6
          30695 => x"81", -- $077e7
          30696 => x"81", -- $077e8
          30697 => x"81", -- $077e9
          30698 => x"81", -- $077ea
          30699 => x"81", -- $077eb
          30700 => x"81", -- $077ec
          30701 => x"80", -- $077ed
          30702 => x"80", -- $077ee
          30703 => x"80", -- $077ef
          30704 => x"80", -- $077f0
          30705 => x"80", -- $077f1
          30706 => x"80", -- $077f2
          30707 => x"80", -- $077f3
          30708 => x"80", -- $077f4
          30709 => x"80", -- $077f5
          30710 => x"80", -- $077f6
          30711 => x"80", -- $077f7
          30712 => x"80", -- $077f8
          30713 => x"80", -- $077f9
          30714 => x"80", -- $077fa
          30715 => x"80", -- $077fb
          30716 => x"80", -- $077fc
          30717 => x"80", -- $077fd
          30718 => x"80", -- $077fe
          30719 => x"80", -- $077ff
          30720 => x"81", -- $07800
          30721 => x"81", -- $07801
          30722 => x"81", -- $07802
          30723 => x"81", -- $07803
          30724 => x"81", -- $07804
          30725 => x"82", -- $07805
          30726 => x"82", -- $07806
          30727 => x"82", -- $07807
          30728 => x"82", -- $07808
          30729 => x"82", -- $07809
          30730 => x"82", -- $0780a
          30731 => x"82", -- $0780b
          30732 => x"82", -- $0780c
          30733 => x"82", -- $0780d
          30734 => x"82", -- $0780e
          30735 => x"82", -- $0780f
          30736 => x"82", -- $07810
          30737 => x"82", -- $07811
          30738 => x"82", -- $07812
          30739 => x"82", -- $07813
          30740 => x"82", -- $07814
          30741 => x"81", -- $07815
          30742 => x"81", -- $07816
          30743 => x"81", -- $07817
          30744 => x"81", -- $07818
          30745 => x"81", -- $07819
          30746 => x"81", -- $0781a
          30747 => x"81", -- $0781b
          30748 => x"81", -- $0781c
          30749 => x"81", -- $0781d
          30750 => x"81", -- $0781e
          30751 => x"81", -- $0781f
          30752 => x"81", -- $07820
          30753 => x"81", -- $07821
          30754 => x"81", -- $07822
          30755 => x"81", -- $07823
          30756 => x"81", -- $07824
          30757 => x"82", -- $07825
          30758 => x"82", -- $07826
          30759 => x"82", -- $07827
          30760 => x"82", -- $07828
          30761 => x"82", -- $07829
          30762 => x"82", -- $0782a
          30763 => x"83", -- $0782b
          30764 => x"83", -- $0782c
          30765 => x"83", -- $0782d
          30766 => x"83", -- $0782e
          30767 => x"83", -- $0782f
          30768 => x"83", -- $07830
          30769 => x"83", -- $07831
          30770 => x"83", -- $07832
          30771 => x"82", -- $07833
          30772 => x"82", -- $07834
          30773 => x"82", -- $07835
          30774 => x"82", -- $07836
          30775 => x"82", -- $07837
          30776 => x"81", -- $07838
          30777 => x"81", -- $07839
          30778 => x"81", -- $0783a
          30779 => x"81", -- $0783b
          30780 => x"81", -- $0783c
          30781 => x"81", -- $0783d
          30782 => x"81", -- $0783e
          30783 => x"81", -- $0783f
          30784 => x"81", -- $07840
          30785 => x"81", -- $07841
          30786 => x"81", -- $07842
          30787 => x"81", -- $07843
          30788 => x"81", -- $07844
          30789 => x"81", -- $07845
          30790 => x"81", -- $07846
          30791 => x"81", -- $07847
          30792 => x"81", -- $07848
          30793 => x"81", -- $07849
          30794 => x"82", -- $0784a
          30795 => x"82", -- $0784b
          30796 => x"82", -- $0784c
          30797 => x"82", -- $0784d
          30798 => x"82", -- $0784e
          30799 => x"82", -- $0784f
          30800 => x"82", -- $07850
          30801 => x"82", -- $07851
          30802 => x"82", -- $07852
          30803 => x"82", -- $07853
          30804 => x"82", -- $07854
          30805 => x"82", -- $07855
          30806 => x"82", -- $07856
          30807 => x"82", -- $07857
          30808 => x"82", -- $07858
          30809 => x"82", -- $07859
          30810 => x"82", -- $0785a
          30811 => x"81", -- $0785b
          30812 => x"81", -- $0785c
          30813 => x"81", -- $0785d
          30814 => x"81", -- $0785e
          30815 => x"81", -- $0785f
          30816 => x"80", -- $07860
          30817 => x"81", -- $07861
          30818 => x"80", -- $07862
          30819 => x"80", -- $07863
          30820 => x"80", -- $07864
          30821 => x"81", -- $07865
          30822 => x"81", -- $07866
          30823 => x"80", -- $07867
          30824 => x"81", -- $07868
          30825 => x"81", -- $07869
          30826 => x"81", -- $0786a
          30827 => x"81", -- $0786b
          30828 => x"81", -- $0786c
          30829 => x"81", -- $0786d
          30830 => x"81", -- $0786e
          30831 => x"82", -- $0786f
          30832 => x"82", -- $07870
          30833 => x"82", -- $07871
          30834 => x"82", -- $07872
          30835 => x"82", -- $07873
          30836 => x"82", -- $07874
          30837 => x"82", -- $07875
          30838 => x"83", -- $07876
          30839 => x"83", -- $07877
          30840 => x"82", -- $07878
          30841 => x"82", -- $07879
          30842 => x"82", -- $0787a
          30843 => x"82", -- $0787b
          30844 => x"82", -- $0787c
          30845 => x"82", -- $0787d
          30846 => x"82", -- $0787e
          30847 => x"82", -- $0787f
          30848 => x"82", -- $07880
          30849 => x"81", -- $07881
          30850 => x"81", -- $07882
          30851 => x"81", -- $07883
          30852 => x"81", -- $07884
          30853 => x"81", -- $07885
          30854 => x"81", -- $07886
          30855 => x"81", -- $07887
          30856 => x"81", -- $07888
          30857 => x"81", -- $07889
          30858 => x"81", -- $0788a
          30859 => x"81", -- $0788b
          30860 => x"81", -- $0788c
          30861 => x"81", -- $0788d
          30862 => x"81", -- $0788e
          30863 => x"81", -- $0788f
          30864 => x"82", -- $07890
          30865 => x"82", -- $07891
          30866 => x"82", -- $07892
          30867 => x"82", -- $07893
          30868 => x"82", -- $07894
          30869 => x"82", -- $07895
          30870 => x"83", -- $07896
          30871 => x"83", -- $07897
          30872 => x"83", -- $07898
          30873 => x"83", -- $07899
          30874 => x"83", -- $0789a
          30875 => x"83", -- $0789b
          30876 => x"83", -- $0789c
          30877 => x"83", -- $0789d
          30878 => x"83", -- $0789e
          30879 => x"83", -- $0789f
          30880 => x"82", -- $078a0
          30881 => x"82", -- $078a1
          30882 => x"82", -- $078a2
          30883 => x"82", -- $078a3
          30884 => x"82", -- $078a4
          30885 => x"82", -- $078a5
          30886 => x"82", -- $078a6
          30887 => x"82", -- $078a7
          30888 => x"81", -- $078a8
          30889 => x"81", -- $078a9
          30890 => x"81", -- $078aa
          30891 => x"81", -- $078ab
          30892 => x"81", -- $078ac
          30893 => x"81", -- $078ad
          30894 => x"81", -- $078ae
          30895 => x"81", -- $078af
          30896 => x"81", -- $078b0
          30897 => x"81", -- $078b1
          30898 => x"81", -- $078b2
          30899 => x"82", -- $078b3
          30900 => x"82", -- $078b4
          30901 => x"82", -- $078b5
          30902 => x"82", -- $078b6
          30903 => x"82", -- $078b7
          30904 => x"83", -- $078b8
          30905 => x"83", -- $078b9
          30906 => x"83", -- $078ba
          30907 => x"83", -- $078bb
          30908 => x"83", -- $078bc
          30909 => x"83", -- $078bd
          30910 => x"83", -- $078be
          30911 => x"83", -- $078bf
          30912 => x"83", -- $078c0
          30913 => x"83", -- $078c1
          30914 => x"83", -- $078c2
          30915 => x"83", -- $078c3
          30916 => x"82", -- $078c4
          30917 => x"82", -- $078c5
          30918 => x"82", -- $078c6
          30919 => x"82", -- $078c7
          30920 => x"82", -- $078c8
          30921 => x"81", -- $078c9
          30922 => x"81", -- $078ca
          30923 => x"81", -- $078cb
          30924 => x"81", -- $078cc
          30925 => x"81", -- $078cd
          30926 => x"81", -- $078ce
          30927 => x"81", -- $078cf
          30928 => x"81", -- $078d0
          30929 => x"81", -- $078d1
          30930 => x"81", -- $078d2
          30931 => x"81", -- $078d3
          30932 => x"81", -- $078d4
          30933 => x"81", -- $078d5
          30934 => x"81", -- $078d6
          30935 => x"82", -- $078d7
          30936 => x"82", -- $078d8
          30937 => x"82", -- $078d9
          30938 => x"82", -- $078da
          30939 => x"82", -- $078db
          30940 => x"83", -- $078dc
          30941 => x"83", -- $078dd
          30942 => x"83", -- $078de
          30943 => x"83", -- $078df
          30944 => x"83", -- $078e0
          30945 => x"83", -- $078e1
          30946 => x"83", -- $078e2
          30947 => x"83", -- $078e3
          30948 => x"83", -- $078e4
          30949 => x"83", -- $078e5
          30950 => x"82", -- $078e6
          30951 => x"82", -- $078e7
          30952 => x"82", -- $078e8
          30953 => x"82", -- $078e9
          30954 => x"81", -- $078ea
          30955 => x"81", -- $078eb
          30956 => x"81", -- $078ec
          30957 => x"81", -- $078ed
          30958 => x"81", -- $078ee
          30959 => x"81", -- $078ef
          30960 => x"80", -- $078f0
          30961 => x"80", -- $078f1
          30962 => x"81", -- $078f2
          30963 => x"81", -- $078f3
          30964 => x"80", -- $078f4
          30965 => x"81", -- $078f5
          30966 => x"81", -- $078f6
          30967 => x"81", -- $078f7
          30968 => x"81", -- $078f8
          30969 => x"81", -- $078f9
          30970 => x"81", -- $078fa
          30971 => x"81", -- $078fb
          30972 => x"81", -- $078fc
          30973 => x"82", -- $078fd
          30974 => x"82", -- $078fe
          30975 => x"82", -- $078ff
          30976 => x"82", -- $07900
          30977 => x"82", -- $07901
          30978 => x"82", -- $07902
          30979 => x"82", -- $07903
          30980 => x"83", -- $07904
          30981 => x"82", -- $07905
          30982 => x"82", -- $07906
          30983 => x"82", -- $07907
          30984 => x"82", -- $07908
          30985 => x"82", -- $07909
          30986 => x"81", -- $0790a
          30987 => x"81", -- $0790b
          30988 => x"81", -- $0790c
          30989 => x"81", -- $0790d
          30990 => x"81", -- $0790e
          30991 => x"81", -- $0790f
          30992 => x"81", -- $07910
          30993 => x"80", -- $07911
          30994 => x"80", -- $07912
          30995 => x"80", -- $07913
          30996 => x"80", -- $07914
          30997 => x"80", -- $07915
          30998 => x"80", -- $07916
          30999 => x"80", -- $07917
          31000 => x"80", -- $07918
          31001 => x"80", -- $07919
          31002 => x"80", -- $0791a
          31003 => x"80", -- $0791b
          31004 => x"80", -- $0791c
          31005 => x"80", -- $0791d
          31006 => x"81", -- $0791e
          31007 => x"81", -- $0791f
          31008 => x"81", -- $07920
          31009 => x"81", -- $07921
          31010 => x"81", -- $07922
          31011 => x"81", -- $07923
          31012 => x"81", -- $07924
          31013 => x"81", -- $07925
          31014 => x"81", -- $07926
          31015 => x"81", -- $07927
          31016 => x"81", -- $07928
          31017 => x"81", -- $07929
          31018 => x"81", -- $0792a
          31019 => x"81", -- $0792b
          31020 => x"81", -- $0792c
          31021 => x"81", -- $0792d
          31022 => x"80", -- $0792e
          31023 => x"80", -- $0792f
          31024 => x"80", -- $07930
          31025 => x"80", -- $07931
          31026 => x"80", -- $07932
          31027 => x"80", -- $07933
          31028 => x"80", -- $07934
          31029 => x"80", -- $07935
          31030 => x"80", -- $07936
          31031 => x"80", -- $07937
          31032 => x"80", -- $07938
          31033 => x"80", -- $07939
          31034 => x"80", -- $0793a
          31035 => x"80", -- $0793b
          31036 => x"80", -- $0793c
          31037 => x"80", -- $0793d
          31038 => x"80", -- $0793e
          31039 => x"80", -- $0793f
          31040 => x"80", -- $07940
          31041 => x"80", -- $07941
          31042 => x"80", -- $07942
          31043 => x"80", -- $07943
          31044 => x"80", -- $07944
          31045 => x"80", -- $07945
          31046 => x"80", -- $07946
          31047 => x"80", -- $07947
          31048 => x"80", -- $07948
          31049 => x"80", -- $07949
          31050 => x"80", -- $0794a
          31051 => x"80", -- $0794b
          31052 => x"80", -- $0794c
          31053 => x"80", -- $0794d
          31054 => x"80", -- $0794e
          31055 => x"80", -- $0794f
          31056 => x"80", -- $07950
          31057 => x"80", -- $07951
          31058 => x"80", -- $07952
          31059 => x"80", -- $07953
          31060 => x"80", -- $07954
          31061 => x"7f", -- $07955
          31062 => x"7f", -- $07956
          31063 => x"7f", -- $07957
          31064 => x"7f", -- $07958
          31065 => x"7f", -- $07959
          31066 => x"7f", -- $0795a
          31067 => x"7f", -- $0795b
          31068 => x"7f", -- $0795c
          31069 => x"7f", -- $0795d
          31070 => x"7f", -- $0795e
          31071 => x"7f", -- $0795f
          31072 => x"7f", -- $07960
          31073 => x"80", -- $07961
          31074 => x"80", -- $07962
          31075 => x"7f", -- $07963
          31076 => x"80", -- $07964
          31077 => x"80", -- $07965
          31078 => x"80", -- $07966
          31079 => x"80", -- $07967
          31080 => x"80", -- $07968
          31081 => x"80", -- $07969
          31082 => x"80", -- $0796a
          31083 => x"80", -- $0796b
          31084 => x"80", -- $0796c
          31085 => x"80", -- $0796d
          31086 => x"80", -- $0796e
          31087 => x"80", -- $0796f
          31088 => x"80", -- $07970
          31089 => x"80", -- $07971
          31090 => x"80", -- $07972
          31091 => x"80", -- $07973
          31092 => x"7f", -- $07974
          31093 => x"80", -- $07975
          31094 => x"7f", -- $07976
          31095 => x"7f", -- $07977
          31096 => x"7f", -- $07978
          31097 => x"7f", -- $07979
          31098 => x"7f", -- $0797a
          31099 => x"7f", -- $0797b
          31100 => x"7f", -- $0797c
          31101 => x"7f", -- $0797d
          31102 => x"7f", -- $0797e
          31103 => x"7f", -- $0797f
          31104 => x"7f", -- $07980
          31105 => x"7f", -- $07981
          31106 => x"7f", -- $07982
          31107 => x"7f", -- $07983
          31108 => x"7f", -- $07984
          31109 => x"7f", -- $07985
          31110 => x"80", -- $07986
          31111 => x"80", -- $07987
          31112 => x"80", -- $07988
          31113 => x"80", -- $07989
          31114 => x"80", -- $0798a
          31115 => x"80", -- $0798b
          31116 => x"80", -- $0798c
          31117 => x"80", -- $0798d
          31118 => x"80", -- $0798e
          31119 => x"80", -- $0798f
          31120 => x"80", -- $07990
          31121 => x"80", -- $07991
          31122 => x"80", -- $07992
          31123 => x"7f", -- $07993
          31124 => x"80", -- $07994
          31125 => x"7f", -- $07995
          31126 => x"7f", -- $07996
          31127 => x"7f", -- $07997
          31128 => x"7f", -- $07998
          31129 => x"7f", -- $07999
          31130 => x"7f", -- $0799a
          31131 => x"7f", -- $0799b
          31132 => x"7f", -- $0799c
          31133 => x"7f", -- $0799d
          31134 => x"7f", -- $0799e
          31135 => x"7f", -- $0799f
          31136 => x"7f", -- $079a0
          31137 => x"7f", -- $079a1
          31138 => x"7f", -- $079a2
          31139 => x"7f", -- $079a3
          31140 => x"7f", -- $079a4
          31141 => x"7f", -- $079a5
          31142 => x"7f", -- $079a6
          31143 => x"7f", -- $079a7
          31144 => x"7f", -- $079a8
          31145 => x"7f", -- $079a9
          31146 => x"7f", -- $079aa
          31147 => x"7f", -- $079ab
          31148 => x"7f", -- $079ac
          31149 => x"7f", -- $079ad
          31150 => x"7f", -- $079ae
          31151 => x"7f", -- $079af
          31152 => x"7f", -- $079b0
          31153 => x"7f", -- $079b1
          31154 => x"7f", -- $079b2
          31155 => x"7f", -- $079b3
          31156 => x"7f", -- $079b4
          31157 => x"7f", -- $079b5
          31158 => x"7f", -- $079b6
          31159 => x"7f", -- $079b7
          31160 => x"7f", -- $079b8
          31161 => x"7f", -- $079b9
          31162 => x"7f", -- $079ba
          31163 => x"7f", -- $079bb
          31164 => x"7f", -- $079bc
          31165 => x"7f", -- $079bd
          31166 => x"7f", -- $079be
          31167 => x"7f", -- $079bf
          31168 => x"7f", -- $079c0
          31169 => x"7f", -- $079c1
          31170 => x"7f", -- $079c2
          31171 => x"7f", -- $079c3
          31172 => x"7f", -- $079c4
          31173 => x"7f", -- $079c5
          31174 => x"80", -- $079c6
          31175 => x"80", -- $079c7
          31176 => x"80", -- $079c8
          31177 => x"80", -- $079c9
          31178 => x"80", -- $079ca
          31179 => x"7f", -- $079cb
          31180 => x"7f", -- $079cc
          31181 => x"7f", -- $079cd
          31182 => x"7f", -- $079ce
          31183 => x"7f", -- $079cf
          31184 => x"7f", -- $079d0
          31185 => x"7f", -- $079d1
          31186 => x"7f", -- $079d2
          31187 => x"7f", -- $079d3
          31188 => x"7f", -- $079d4
          31189 => x"7f", -- $079d5
          31190 => x"7f", -- $079d6
          31191 => x"7f", -- $079d7
          31192 => x"7f", -- $079d8
          31193 => x"7f", -- $079d9
          31194 => x"7f", -- $079da
          31195 => x"7f", -- $079db
          31196 => x"7f", -- $079dc
          31197 => x"7f", -- $079dd
          31198 => x"7f", -- $079de
          31199 => x"7f", -- $079df
          31200 => x"7f", -- $079e0
          31201 => x"7f", -- $079e1
          31202 => x"7f", -- $079e2
          31203 => x"7f", -- $079e3
          31204 => x"7f", -- $079e4
          31205 => x"7f", -- $079e5
          31206 => x"7f", -- $079e6
          31207 => x"7f", -- $079e7
          31208 => x"7f", -- $079e8
          31209 => x"7f", -- $079e9
          31210 => x"7f", -- $079ea
          31211 => x"7f", -- $079eb
          31212 => x"7f", -- $079ec
          31213 => x"7f", -- $079ed
          31214 => x"7f", -- $079ee
          31215 => x"7e", -- $079ef
          31216 => x"7e", -- $079f0
          31217 => x"7e", -- $079f1
          31218 => x"7e", -- $079f2
          31219 => x"7e", -- $079f3
          31220 => x"7e", -- $079f4
          31221 => x"7e", -- $079f5
          31222 => x"7e", -- $079f6
          31223 => x"7e", -- $079f7
          31224 => x"7e", -- $079f8
          31225 => x"7e", -- $079f9
          31226 => x"7e", -- $079fa
          31227 => x"7e", -- $079fb
          31228 => x"7e", -- $079fc
          31229 => x"7e", -- $079fd
          31230 => x"7e", -- $079fe
          31231 => x"7e", -- $079ff
          31232 => x"7e", -- $07a00
          31233 => x"7e", -- $07a01
          31234 => x"7e", -- $07a02
          31235 => x"7e", -- $07a03
          31236 => x"7e", -- $07a04
          31237 => x"7f", -- $07a05
          31238 => x"7f", -- $07a06
          31239 => x"7e", -- $07a07
          31240 => x"7f", -- $07a08
          31241 => x"7f", -- $07a09
          31242 => x"7f", -- $07a0a
          31243 => x"7e", -- $07a0b
          31244 => x"7e", -- $07a0c
          31245 => x"7e", -- $07a0d
          31246 => x"7e", -- $07a0e
          31247 => x"7e", -- $07a0f
          31248 => x"7e", -- $07a10
          31249 => x"7d", -- $07a11
          31250 => x"7d", -- $07a12
          31251 => x"7d", -- $07a13
          31252 => x"7d", -- $07a14
          31253 => x"7d", -- $07a15
          31254 => x"7c", -- $07a16
          31255 => x"7c", -- $07a17
          31256 => x"7c", -- $07a18
          31257 => x"7c", -- $07a19
          31258 => x"7c", -- $07a1a
          31259 => x"7c", -- $07a1b
          31260 => x"7d", -- $07a1c
          31261 => x"7d", -- $07a1d
          31262 => x"7d", -- $07a1e
          31263 => x"7d", -- $07a1f
          31264 => x"7d", -- $07a20
          31265 => x"7e", -- $07a21
          31266 => x"7e", -- $07a22
          31267 => x"7e", -- $07a23
          31268 => x"7e", -- $07a24
          31269 => x"7e", -- $07a25
          31270 => x"7e", -- $07a26
          31271 => x"7e", -- $07a27
          31272 => x"7e", -- $07a28
          31273 => x"7e", -- $07a29
          31274 => x"7e", -- $07a2a
          31275 => x"7e", -- $07a2b
          31276 => x"7e", -- $07a2c
          31277 => x"7e", -- $07a2d
          31278 => x"7e", -- $07a2e
          31279 => x"7d", -- $07a2f
          31280 => x"7d", -- $07a30
          31281 => x"7d", -- $07a31
          31282 => x"7d", -- $07a32
          31283 => x"7d", -- $07a33
          31284 => x"7c", -- $07a34
          31285 => x"7c", -- $07a35
          31286 => x"7c", -- $07a36
          31287 => x"7c", -- $07a37
          31288 => x"7c", -- $07a38
          31289 => x"7c", -- $07a39
          31290 => x"7c", -- $07a3a
          31291 => x"7c", -- $07a3b
          31292 => x"7c", -- $07a3c
          31293 => x"7c", -- $07a3d
          31294 => x"7d", -- $07a3e
          31295 => x"7d", -- $07a3f
          31296 => x"7d", -- $07a40
          31297 => x"7d", -- $07a41
          31298 => x"7d", -- $07a42
          31299 => x"7e", -- $07a43
          31300 => x"7e", -- $07a44
          31301 => x"7e", -- $07a45
          31302 => x"7e", -- $07a46
          31303 => x"7e", -- $07a47
          31304 => x"7e", -- $07a48
          31305 => x"7f", -- $07a49
          31306 => x"7f", -- $07a4a
          31307 => x"7e", -- $07a4b
          31308 => x"7e", -- $07a4c
          31309 => x"7e", -- $07a4d
          31310 => x"7e", -- $07a4e
          31311 => x"7e", -- $07a4f
          31312 => x"7e", -- $07a50
          31313 => x"7d", -- $07a51
          31314 => x"7d", -- $07a52
          31315 => x"7d", -- $07a53
          31316 => x"7d", -- $07a54
          31317 => x"7d", -- $07a55
          31318 => x"7d", -- $07a56
          31319 => x"7d", -- $07a57
          31320 => x"7c", -- $07a58
          31321 => x"7d", -- $07a59
          31322 => x"7d", -- $07a5a
          31323 => x"7d", -- $07a5b
          31324 => x"7d", -- $07a5c
          31325 => x"7d", -- $07a5d
          31326 => x"7d", -- $07a5e
          31327 => x"7d", -- $07a5f
          31328 => x"7e", -- $07a60
          31329 => x"7e", -- $07a61
          31330 => x"7e", -- $07a62
          31331 => x"7e", -- $07a63
          31332 => x"7f", -- $07a64
          31333 => x"7f", -- $07a65
          31334 => x"7f", -- $07a66
          31335 => x"7f", -- $07a67
          31336 => x"7f", -- $07a68
          31337 => x"80", -- $07a69
          31338 => x"80", -- $07a6a
          31339 => x"80", -- $07a6b
          31340 => x"7f", -- $07a6c
          31341 => x"7f", -- $07a6d
          31342 => x"7f", -- $07a6e
          31343 => x"7f", -- $07a6f
          31344 => x"7f", -- $07a70
          31345 => x"7f", -- $07a71
          31346 => x"7f", -- $07a72
          31347 => x"7e", -- $07a73
          31348 => x"7e", -- $07a74
          31349 => x"7e", -- $07a75
          31350 => x"7e", -- $07a76
          31351 => x"7e", -- $07a77
          31352 => x"7e", -- $07a78
          31353 => x"7e", -- $07a79
          31354 => x"7e", -- $07a7a
          31355 => x"7e", -- $07a7b
          31356 => x"7e", -- $07a7c
          31357 => x"7e", -- $07a7d
          31358 => x"7e", -- $07a7e
          31359 => x"7e", -- $07a7f
          31360 => x"7f", -- $07a80
          31361 => x"7f", -- $07a81
          31362 => x"7f", -- $07a82
          31363 => x"7f", -- $07a83
          31364 => x"80", -- $07a84
          31365 => x"80", -- $07a85
          31366 => x"80", -- $07a86
          31367 => x"80", -- $07a87
          31368 => x"80", -- $07a88
          31369 => x"80", -- $07a89
          31370 => x"80", -- $07a8a
          31371 => x"80", -- $07a8b
          31372 => x"80", -- $07a8c
          31373 => x"80", -- $07a8d
          31374 => x"80", -- $07a8e
          31375 => x"80", -- $07a8f
          31376 => x"80", -- $07a90
          31377 => x"80", -- $07a91
          31378 => x"80", -- $07a92
          31379 => x"80", -- $07a93
          31380 => x"80", -- $07a94
          31381 => x"80", -- $07a95
          31382 => x"7f", -- $07a96
          31383 => x"7f", -- $07a97
          31384 => x"7f", -- $07a98
          31385 => x"7f", -- $07a99
          31386 => x"7f", -- $07a9a
          31387 => x"7f", -- $07a9b
          31388 => x"7f", -- $07a9c
          31389 => x"7f", -- $07a9d
          31390 => x"7f", -- $07a9e
          31391 => x"80", -- $07a9f
          31392 => x"80", -- $07aa0
          31393 => x"80", -- $07aa1
          31394 => x"80", -- $07aa2
          31395 => x"80", -- $07aa3
          31396 => x"80", -- $07aa4
          31397 => x"80", -- $07aa5
          31398 => x"80", -- $07aa6
          31399 => x"80", -- $07aa7
          31400 => x"80", -- $07aa8
          31401 => x"80", -- $07aa9
          31402 => x"80", -- $07aaa
          31403 => x"80", -- $07aab
          31404 => x"80", -- $07aac
          31405 => x"80", -- $07aad
          31406 => x"80", -- $07aae
          31407 => x"80", -- $07aaf
          31408 => x"80", -- $07ab0
          31409 => x"80", -- $07ab1
          31410 => x"80", -- $07ab2
          31411 => x"80", -- $07ab3
          31412 => x"80", -- $07ab4
          31413 => x"80", -- $07ab5
          31414 => x"80", -- $07ab6
          31415 => x"80", -- $07ab7
          31416 => x"80", -- $07ab8
          31417 => x"80", -- $07ab9
          31418 => x"80", -- $07aba
          31419 => x"80", -- $07abb
          31420 => x"80", -- $07abc
          31421 => x"80", -- $07abd
          31422 => x"80", -- $07abe
          31423 => x"80", -- $07abf
          31424 => x"80", -- $07ac0
          31425 => x"80", -- $07ac1
          31426 => x"80", -- $07ac2
          31427 => x"80", -- $07ac3
          31428 => x"80", -- $07ac4
          31429 => x"80", -- $07ac5
          31430 => x"80", -- $07ac6
          31431 => x"80", -- $07ac7
          31432 => x"80", -- $07ac8
          31433 => x"81", -- $07ac9
          31434 => x"81", -- $07aca
          31435 => x"81", -- $07acb
          31436 => x"81", -- $07acc
          31437 => x"81", -- $07acd
          31438 => x"81", -- $07ace
          31439 => x"81", -- $07acf
          31440 => x"80", -- $07ad0
          31441 => x"80", -- $07ad1
          31442 => x"80", -- $07ad2
          31443 => x"80", -- $07ad3
          31444 => x"80", -- $07ad4
          31445 => x"80", -- $07ad5
          31446 => x"80", -- $07ad6
          31447 => x"80", -- $07ad7
          31448 => x"80", -- $07ad8
          31449 => x"80", -- $07ad9
          31450 => x"80", -- $07ada
          31451 => x"80", -- $07adb
          31452 => x"80", -- $07adc
          31453 => x"80", -- $07add
          31454 => x"80", -- $07ade
          31455 => x"80", -- $07adf
          31456 => x"80", -- $07ae0
          31457 => x"80", -- $07ae1
          31458 => x"80", -- $07ae2
          31459 => x"80", -- $07ae3
          31460 => x"80", -- $07ae4
          31461 => x"80", -- $07ae5
          31462 => x"80", -- $07ae6
          31463 => x"80", -- $07ae7
          31464 => x"80", -- $07ae8
          31465 => x"80", -- $07ae9
          31466 => x"80", -- $07aea
          31467 => x"80", -- $07aeb
          31468 => x"80", -- $07aec
          31469 => x"81", -- $07aed
          31470 => x"81", -- $07aee
          31471 => x"81", -- $07aef
          31472 => x"80", -- $07af0
          31473 => x"80", -- $07af1
          31474 => x"80", -- $07af2
          31475 => x"80", -- $07af3
          31476 => x"80", -- $07af4
          31477 => x"80", -- $07af5
          31478 => x"80", -- $07af6
          31479 => x"80", -- $07af7
          31480 => x"80", -- $07af8
          31481 => x"80", -- $07af9
          31482 => x"80", -- $07afa
          31483 => x"80", -- $07afb
          31484 => x"80", -- $07afc
          31485 => x"80", -- $07afd
          31486 => x"80", -- $07afe
          31487 => x"80", -- $07aff
          31488 => x"80", -- $07b00
          31489 => x"80", -- $07b01
          31490 => x"80", -- $07b02
          31491 => x"80", -- $07b03
          31492 => x"80", -- $07b04
          31493 => x"80", -- $07b05
          31494 => x"80", -- $07b06
          31495 => x"80", -- $07b07
          31496 => x"80", -- $07b08
          31497 => x"81", -- $07b09
          31498 => x"81", -- $07b0a
          31499 => x"81", -- $07b0b
          31500 => x"81", -- $07b0c
          31501 => x"81", -- $07b0d
          31502 => x"81", -- $07b0e
          31503 => x"81", -- $07b0f
          31504 => x"81", -- $07b10
          31505 => x"81", -- $07b11
          31506 => x"80", -- $07b12
          31507 => x"80", -- $07b13
          31508 => x"80", -- $07b14
          31509 => x"80", -- $07b15
          31510 => x"80", -- $07b16
          31511 => x"80", -- $07b17
          31512 => x"80", -- $07b18
          31513 => x"80", -- $07b19
          31514 => x"80", -- $07b1a
          31515 => x"80", -- $07b1b
          31516 => x"80", -- $07b1c
          31517 => x"80", -- $07b1d
          31518 => x"80", -- $07b1e
          31519 => x"81", -- $07b1f
          31520 => x"81", -- $07b20
          31521 => x"81", -- $07b21
          31522 => x"81", -- $07b22
          31523 => x"81", -- $07b23
          31524 => x"81", -- $07b24
          31525 => x"81", -- $07b25
          31526 => x"81", -- $07b26
          31527 => x"81", -- $07b27
          31528 => x"81", -- $07b28
          31529 => x"81", -- $07b29
          31530 => x"81", -- $07b2a
          31531 => x"81", -- $07b2b
          31532 => x"81", -- $07b2c
          31533 => x"81", -- $07b2d
          31534 => x"81", -- $07b2e
          31535 => x"81", -- $07b2f
          31536 => x"81", -- $07b30
          31537 => x"81", -- $07b31
          31538 => x"81", -- $07b32
          31539 => x"81", -- $07b33
          31540 => x"81", -- $07b34
          31541 => x"81", -- $07b35
          31542 => x"81", -- $07b36
          31543 => x"80", -- $07b37
          31544 => x"80", -- $07b38
          31545 => x"80", -- $07b39
          31546 => x"80", -- $07b3a
          31547 => x"81", -- $07b3b
          31548 => x"81", -- $07b3c
          31549 => x"81", -- $07b3d
          31550 => x"81", -- $07b3e
          31551 => x"81", -- $07b3f
          31552 => x"81", -- $07b40
          31553 => x"82", -- $07b41
          31554 => x"82", -- $07b42
          31555 => x"82", -- $07b43
          31556 => x"82", -- $07b44
          31557 => x"82", -- $07b45
          31558 => x"81", -- $07b46
          31559 => x"82", -- $07b47
          31560 => x"82", -- $07b48
          31561 => x"82", -- $07b49
          31562 => x"82", -- $07b4a
          31563 => x"82", -- $07b4b
          31564 => x"82", -- $07b4c
          31565 => x"82", -- $07b4d
          31566 => x"82", -- $07b4e
          31567 => x"81", -- $07b4f
          31568 => x"81", -- $07b50
          31569 => x"81", -- $07b51
          31570 => x"81", -- $07b52
          31571 => x"81", -- $07b53
          31572 => x"81", -- $07b54
          31573 => x"81", -- $07b55
          31574 => x"81", -- $07b56
          31575 => x"81", -- $07b57
          31576 => x"81", -- $07b58
          31577 => x"81", -- $07b59
          31578 => x"81", -- $07b5a
          31579 => x"81", -- $07b5b
          31580 => x"81", -- $07b5c
          31581 => x"81", -- $07b5d
          31582 => x"81", -- $07b5e
          31583 => x"81", -- $07b5f
          31584 => x"82", -- $07b60
          31585 => x"82", -- $07b61
          31586 => x"82", -- $07b62
          31587 => x"82", -- $07b63
          31588 => x"82", -- $07b64
          31589 => x"82", -- $07b65
          31590 => x"82", -- $07b66
          31591 => x"82", -- $07b67
          31592 => x"82", -- $07b68
          31593 => x"82", -- $07b69
          31594 => x"82", -- $07b6a
          31595 => x"82", -- $07b6b
          31596 => x"82", -- $07b6c
          31597 => x"82", -- $07b6d
          31598 => x"82", -- $07b6e
          31599 => x"82", -- $07b6f
          31600 => x"82", -- $07b70
          31601 => x"82", -- $07b71
          31602 => x"82", -- $07b72
          31603 => x"81", -- $07b73
          31604 => x"81", -- $07b74
          31605 => x"81", -- $07b75
          31606 => x"81", -- $07b76
          31607 => x"81", -- $07b77
          31608 => x"81", -- $07b78
          31609 => x"81", -- $07b79
          31610 => x"81", -- $07b7a
          31611 => x"81", -- $07b7b
          31612 => x"81", -- $07b7c
          31613 => x"81", -- $07b7d
          31614 => x"82", -- $07b7e
          31615 => x"82", -- $07b7f
          31616 => x"82", -- $07b80
          31617 => x"82", -- $07b81
          31618 => x"82", -- $07b82
          31619 => x"83", -- $07b83
          31620 => x"83", -- $07b84
          31621 => x"83", -- $07b85
          31622 => x"83", -- $07b86
          31623 => x"83", -- $07b87
          31624 => x"83", -- $07b88
          31625 => x"83", -- $07b89
          31626 => x"83", -- $07b8a
          31627 => x"83", -- $07b8b
          31628 => x"83", -- $07b8c
          31629 => x"83", -- $07b8d
          31630 => x"83", -- $07b8e
          31631 => x"83", -- $07b8f
          31632 => x"83", -- $07b90
          31633 => x"82", -- $07b91
          31634 => x"82", -- $07b92
          31635 => x"82", -- $07b93
          31636 => x"82", -- $07b94
          31637 => x"82", -- $07b95
          31638 => x"82", -- $07b96
          31639 => x"81", -- $07b97
          31640 => x"81", -- $07b98
          31641 => x"81", -- $07b99
          31642 => x"81", -- $07b9a
          31643 => x"81", -- $07b9b
          31644 => x"81", -- $07b9c
          31645 => x"82", -- $07b9d
          31646 => x"82", -- $07b9e
          31647 => x"82", -- $07b9f
          31648 => x"82", -- $07ba0
          31649 => x"82", -- $07ba1
          31650 => x"82", -- $07ba2
          31651 => x"82", -- $07ba3
          31652 => x"83", -- $07ba4
          31653 => x"83", -- $07ba5
          31654 => x"83", -- $07ba6
          31655 => x"83", -- $07ba7
          31656 => x"83", -- $07ba8
          31657 => x"83", -- $07ba9
          31658 => x"83", -- $07baa
          31659 => x"83", -- $07bab
          31660 => x"83", -- $07bac
          31661 => x"83", -- $07bad
          31662 => x"83", -- $07bae
          31663 => x"82", -- $07baf
          31664 => x"82", -- $07bb0
          31665 => x"82", -- $07bb1
          31666 => x"82", -- $07bb2
          31667 => x"82", -- $07bb3
          31668 => x"82", -- $07bb4
          31669 => x"82", -- $07bb5
          31670 => x"81", -- $07bb6
          31671 => x"81", -- $07bb7
          31672 => x"81", -- $07bb8
          31673 => x"81", -- $07bb9
          31674 => x"81", -- $07bba
          31675 => x"81", -- $07bbb
          31676 => x"81", -- $07bbc
          31677 => x"81", -- $07bbd
          31678 => x"81", -- $07bbe
          31679 => x"81", -- $07bbf
          31680 => x"81", -- $07bc0
          31681 => x"82", -- $07bc1
          31682 => x"82", -- $07bc2
          31683 => x"82", -- $07bc3
          31684 => x"82", -- $07bc4
          31685 => x"82", -- $07bc5
          31686 => x"82", -- $07bc6
          31687 => x"82", -- $07bc7
          31688 => x"82", -- $07bc8
          31689 => x"82", -- $07bc9
          31690 => x"82", -- $07bca
          31691 => x"82", -- $07bcb
          31692 => x"82", -- $07bcc
          31693 => x"82", -- $07bcd
          31694 => x"82", -- $07bce
          31695 => x"82", -- $07bcf
          31696 => x"82", -- $07bd0
          31697 => x"82", -- $07bd1
          31698 => x"81", -- $07bd2
          31699 => x"81", -- $07bd3
          31700 => x"81", -- $07bd4
          31701 => x"81", -- $07bd5
          31702 => x"81", -- $07bd6
          31703 => x"81", -- $07bd7
          31704 => x"81", -- $07bd8
          31705 => x"80", -- $07bd9
          31706 => x"80", -- $07bda
          31707 => x"80", -- $07bdb
          31708 => x"80", -- $07bdc
          31709 => x"81", -- $07bdd
          31710 => x"81", -- $07bde
          31711 => x"80", -- $07bdf
          31712 => x"80", -- $07be0
          31713 => x"81", -- $07be1
          31714 => x"80", -- $07be2
          31715 => x"81", -- $07be3
          31716 => x"81", -- $07be4
          31717 => x"81", -- $07be5
          31718 => x"81", -- $07be6
          31719 => x"81", -- $07be7
          31720 => x"81", -- $07be8
          31721 => x"81", -- $07be9
          31722 => x"81", -- $07bea
          31723 => x"81", -- $07beb
          31724 => x"81", -- $07bec
          31725 => x"81", -- $07bed
          31726 => x"81", -- $07bee
          31727 => x"81", -- $07bef
          31728 => x"81", -- $07bf0
          31729 => x"81", -- $07bf1
          31730 => x"81", -- $07bf2
          31731 => x"81", -- $07bf3
          31732 => x"81", -- $07bf4
          31733 => x"81", -- $07bf5
          31734 => x"81", -- $07bf6
          31735 => x"80", -- $07bf7
          31736 => x"80", -- $07bf8
          31737 => x"80", -- $07bf9
          31738 => x"80", -- $07bfa
          31739 => x"80", -- $07bfb
          31740 => x"80", -- $07bfc
          31741 => x"80", -- $07bfd
          31742 => x"80", -- $07bfe
          31743 => x"80", -- $07bff
          31744 => x"80", -- $07c00
          31745 => x"80", -- $07c01
          31746 => x"80", -- $07c02
          31747 => x"80", -- $07c03
          31748 => x"80", -- $07c04
          31749 => x"80", -- $07c05
          31750 => x"80", -- $07c06
          31751 => x"80", -- $07c07
          31752 => x"80", -- $07c08
          31753 => x"80", -- $07c09
          31754 => x"80", -- $07c0a
          31755 => x"80", -- $07c0b
          31756 => x"80", -- $07c0c
          31757 => x"80", -- $07c0d
          31758 => x"80", -- $07c0e
          31759 => x"80", -- $07c0f
          31760 => x"80", -- $07c10
          31761 => x"80", -- $07c11
          31762 => x"80", -- $07c12
          31763 => x"80", -- $07c13
          31764 => x"80", -- $07c14
          31765 => x"80", -- $07c15
          31766 => x"80", -- $07c16
          31767 => x"80", -- $07c17
          31768 => x"80", -- $07c18
          31769 => x"80", -- $07c19
          31770 => x"80", -- $07c1a
          31771 => x"80", -- $07c1b
          31772 => x"80", -- $07c1c
          31773 => x"80", -- $07c1d
          31774 => x"80", -- $07c1e
          31775 => x"80", -- $07c1f
          31776 => x"80", -- $07c20
          31777 => x"80", -- $07c21
          31778 => x"80", -- $07c22
          31779 => x"80", -- $07c23
          31780 => x"80", -- $07c24
          31781 => x"80", -- $07c25
          31782 => x"80", -- $07c26
          31783 => x"80", -- $07c27
          31784 => x"80", -- $07c28
          31785 => x"80", -- $07c29
          31786 => x"80", -- $07c2a
          31787 => x"80", -- $07c2b
          31788 => x"80", -- $07c2c
          31789 => x"80", -- $07c2d
          31790 => x"80", -- $07c2e
          31791 => x"80", -- $07c2f
          31792 => x"80", -- $07c30
          31793 => x"80", -- $07c31
          31794 => x"80", -- $07c32
          31795 => x"80", -- $07c33
          31796 => x"80", -- $07c34
          31797 => x"80", -- $07c35
          31798 => x"80", -- $07c36
          31799 => x"80", -- $07c37
          31800 => x"80", -- $07c38
          31801 => x"80", -- $07c39
          31802 => x"80", -- $07c3a
          31803 => x"80", -- $07c3b
          31804 => x"80", -- $07c3c
          31805 => x"80", -- $07c3d
          31806 => x"80", -- $07c3e
          31807 => x"80", -- $07c3f
          31808 => x"80", -- $07c40
          31809 => x"80", -- $07c41
          31810 => x"80", -- $07c42
          31811 => x"80", -- $07c43
          31812 => x"80", -- $07c44
          31813 => x"80", -- $07c45
          31814 => x"80", -- $07c46
          31815 => x"80", -- $07c47
          31816 => x"80", -- $07c48
          31817 => x"80", -- $07c49
          31818 => x"80", -- $07c4a
          31819 => x"80", -- $07c4b
          31820 => x"80", -- $07c4c
          31821 => x"80", -- $07c4d
          31822 => x"80", -- $07c4e
          31823 => x"80", -- $07c4f
          31824 => x"80", -- $07c50
          31825 => x"80", -- $07c51
          31826 => x"80", -- $07c52
          31827 => x"80", -- $07c53
          31828 => x"80", -- $07c54
          31829 => x"80", -- $07c55
          31830 => x"80", -- $07c56
          31831 => x"80", -- $07c57
          31832 => x"80", -- $07c58
          31833 => x"80", -- $07c59
          31834 => x"80", -- $07c5a
          31835 => x"80", -- $07c5b
          31836 => x"80", -- $07c5c
          31837 => x"80", -- $07c5d
          31838 => x"80", -- $07c5e
          31839 => x"80", -- $07c5f
          31840 => x"80", -- $07c60
          31841 => x"80", -- $07c61
          31842 => x"80", -- $07c62
          31843 => x"80", -- $07c63
          31844 => x"80", -- $07c64
          31845 => x"80", -- $07c65
          31846 => x"80", -- $07c66
          31847 => x"80", -- $07c67
          31848 => x"80", -- $07c68
          31849 => x"80", -- $07c69
          31850 => x"80", -- $07c6a
          31851 => x"80", -- $07c6b
          31852 => x"80", -- $07c6c
          31853 => x"80", -- $07c6d
          31854 => x"80", -- $07c6e
          31855 => x"80", -- $07c6f
          31856 => x"80", -- $07c70
          31857 => x"80", -- $07c71
          31858 => x"80", -- $07c72
          31859 => x"7f", -- $07c73
          31860 => x"7f", -- $07c74
          31861 => x"7f", -- $07c75
          31862 => x"7f", -- $07c76
          31863 => x"7f", -- $07c77
          31864 => x"7f", -- $07c78
          31865 => x"7f", -- $07c79
          31866 => x"7f", -- $07c7a
          31867 => x"7f", -- $07c7b
          31868 => x"7f", -- $07c7c
          31869 => x"7f", -- $07c7d
          31870 => x"7f", -- $07c7e
          31871 => x"7f", -- $07c7f
          31872 => x"7f", -- $07c80
          31873 => x"7f", -- $07c81
          31874 => x"7f", -- $07c82
          31875 => x"7f", -- $07c83
          31876 => x"7f", -- $07c84
          31877 => x"7f", -- $07c85
          31878 => x"80", -- $07c86
          31879 => x"7f", -- $07c87
          31880 => x"80", -- $07c88
          31881 => x"7f", -- $07c89
          31882 => x"80", -- $07c8a
          31883 => x"7f", -- $07c8b
          31884 => x"7f", -- $07c8c
          31885 => x"7f", -- $07c8d
          31886 => x"7f", -- $07c8e
          31887 => x"7f", -- $07c8f
          31888 => x"7f", -- $07c90
          31889 => x"7f", -- $07c91
          31890 => x"7f", -- $07c92
          31891 => x"7f", -- $07c93
          31892 => x"7f", -- $07c94
          31893 => x"7e", -- $07c95
          31894 => x"7e", -- $07c96
          31895 => x"7e", -- $07c97
          31896 => x"7e", -- $07c98
          31897 => x"7e", -- $07c99
          31898 => x"7e", -- $07c9a
          31899 => x"7e", -- $07c9b
          31900 => x"7e", -- $07c9c
          31901 => x"7e", -- $07c9d
          31902 => x"7e", -- $07c9e
          31903 => x"7e", -- $07c9f
          31904 => x"7e", -- $07ca0
          31905 => x"7e", -- $07ca1
          31906 => x"7e", -- $07ca2
          31907 => x"7f", -- $07ca3
          31908 => x"7f", -- $07ca4
          31909 => x"7f", -- $07ca5
          31910 => x"7f", -- $07ca6
          31911 => x"7f", -- $07ca7
          31912 => x"7f", -- $07ca8
          31913 => x"7f", -- $07ca9
          31914 => x"80", -- $07caa
          31915 => x"80", -- $07cab
          31916 => x"80", -- $07cac
          31917 => x"80", -- $07cad
          31918 => x"80", -- $07cae
          31919 => x"7f", -- $07caf
          31920 => x"7f", -- $07cb0
          31921 => x"7f", -- $07cb1
          31922 => x"7f", -- $07cb2
          31923 => x"7e", -- $07cb3
          31924 => x"7e", -- $07cb4
          31925 => x"7e", -- $07cb5
          31926 => x"7e", -- $07cb6
          31927 => x"7e", -- $07cb7
          31928 => x"7e", -- $07cb8
          31929 => x"7e", -- $07cb9
          31930 => x"7d", -- $07cba
          31931 => x"7d", -- $07cbb
          31932 => x"7d", -- $07cbc
          31933 => x"7d", -- $07cbd
          31934 => x"7d", -- $07cbe
          31935 => x"7d", -- $07cbf
          31936 => x"7e", -- $07cc0
          31937 => x"7e", -- $07cc1
          31938 => x"7e", -- $07cc2
          31939 => x"7e", -- $07cc3
          31940 => x"7f", -- $07cc4
          31941 => x"7f", -- $07cc5
          31942 => x"7f", -- $07cc6
          31943 => x"7f", -- $07cc7
          31944 => x"7f", -- $07cc8
          31945 => x"80", -- $07cc9
          31946 => x"80", -- $07cca
          31947 => x"80", -- $07ccb
          31948 => x"80", -- $07ccc
          31949 => x"80", -- $07ccd
          31950 => x"80", -- $07cce
          31951 => x"7f", -- $07ccf
          31952 => x"7f", -- $07cd0
          31953 => x"7f", -- $07cd1
          31954 => x"7f", -- $07cd2
          31955 => x"7f", -- $07cd3
          31956 => x"7f", -- $07cd4
          31957 => x"7e", -- $07cd5
          31958 => x"7e", -- $07cd6
          31959 => x"7e", -- $07cd7
          31960 => x"7e", -- $07cd8
          31961 => x"7e", -- $07cd9
          31962 => x"7e", -- $07cda
          31963 => x"7d", -- $07cdb
          31964 => x"7e", -- $07cdc
          31965 => x"7e", -- $07cdd
          31966 => x"7e", -- $07cde
          31967 => x"7e", -- $07cdf
          31968 => x"7e", -- $07ce0
          31969 => x"7e", -- $07ce1
          31970 => x"7e", -- $07ce2
          31971 => x"7f", -- $07ce3
          31972 => x"7f", -- $07ce4
          31973 => x"7f", -- $07ce5
          31974 => x"7f", -- $07ce6
          31975 => x"7f", -- $07ce7
          31976 => x"80", -- $07ce8
          31977 => x"80", -- $07ce9
          31978 => x"80", -- $07cea
          31979 => x"80", -- $07ceb
          31980 => x"80", -- $07cec
          31981 => x"80", -- $07ced
          31982 => x"80", -- $07cee
          31983 => x"80", -- $07cef
          31984 => x"80", -- $07cf0
          31985 => x"7f", -- $07cf1
          31986 => x"7f", -- $07cf2
          31987 => x"7f", -- $07cf3
          31988 => x"7f", -- $07cf4
          31989 => x"7f", -- $07cf5
          31990 => x"7e", -- $07cf6
          31991 => x"7e", -- $07cf7
          31992 => x"7e", -- $07cf8
          31993 => x"7e", -- $07cf9
          31994 => x"7e", -- $07cfa
          31995 => x"7e", -- $07cfb
          31996 => x"7e", -- $07cfc
          31997 => x"7e", -- $07cfd
          31998 => x"7e", -- $07cfe
          31999 => x"7e", -- $07cff
          32000 => x"7e", -- $07d00
          32001 => x"7e", -- $07d01
          32002 => x"7e", -- $07d02
          32003 => x"7e", -- $07d03
          32004 => x"7e", -- $07d04
          32005 => x"7e", -- $07d05
          32006 => x"7f", -- $07d06
          32007 => x"7f", -- $07d07
          32008 => x"7f", -- $07d08
          32009 => x"80", -- $07d09
          32010 => x"80", -- $07d0a
          32011 => x"80", -- $07d0b
          32012 => x"80", -- $07d0c
          32013 => x"80", -- $07d0d
          32014 => x"80", -- $07d0e
          32015 => x"80", -- $07d0f
          32016 => x"80", -- $07d10
          32017 => x"7f", -- $07d11
          32018 => x"7f", -- $07d12
          32019 => x"7f", -- $07d13
          32020 => x"7f", -- $07d14
          32021 => x"7f", -- $07d15
          32022 => x"7f", -- $07d16
          32023 => x"7f", -- $07d17
          32024 => x"7e", -- $07d18
          32025 => x"7e", -- $07d19
          32026 => x"7e", -- $07d1a
          32027 => x"7e", -- $07d1b
          32028 => x"7d", -- $07d1c
          32029 => x"7d", -- $07d1d
          32030 => x"7d", -- $07d1e
          32031 => x"7e", -- $07d1f
          32032 => x"7d", -- $07d20
          32033 => x"7e", -- $07d21
          32034 => x"7e", -- $07d22
          32035 => x"7e", -- $07d23
          32036 => x"7e", -- $07d24
          32037 => x"7e", -- $07d25
          32038 => x"7e", -- $07d26
          32039 => x"7f", -- $07d27
          32040 => x"7f", -- $07d28
          32041 => x"7f", -- $07d29
          32042 => x"7f", -- $07d2a
          32043 => x"7f", -- $07d2b
          32044 => x"80", -- $07d2c
          32045 => x"80", -- $07d2d
          32046 => x"80", -- $07d2e
          32047 => x"80", -- $07d2f
          32048 => x"80", -- $07d30
          32049 => x"80", -- $07d31
          32050 => x"7f", -- $07d32
          32051 => x"7f", -- $07d33
          32052 => x"7f", -- $07d34
          32053 => x"7f", -- $07d35
          32054 => x"7f", -- $07d36
          32055 => x"7f", -- $07d37
          32056 => x"7e", -- $07d38
          32057 => x"7e", -- $07d39
          32058 => x"7e", -- $07d3a
          32059 => x"7e", -- $07d3b
          32060 => x"7e", -- $07d3c
          32061 => x"7e", -- $07d3d
          32062 => x"7e", -- $07d3e
          32063 => x"7e", -- $07d3f
          32064 => x"7e", -- $07d40
          32065 => x"7e", -- $07d41
          32066 => x"7e", -- $07d42
          32067 => x"7e", -- $07d43
          32068 => x"7e", -- $07d44
          32069 => x"7e", -- $07d45
          32070 => x"7f", -- $07d46
          32071 => x"7f", -- $07d47
          32072 => x"7f", -- $07d48
          32073 => x"7f", -- $07d49
          32074 => x"7f", -- $07d4a
          32075 => x"80", -- $07d4b
          32076 => x"80", -- $07d4c
          32077 => x"80", -- $07d4d
          32078 => x"80", -- $07d4e
          32079 => x"80", -- $07d4f
          32080 => x"80", -- $07d50
          32081 => x"80", -- $07d51
          32082 => x"7f", -- $07d52
          32083 => x"80", -- $07d53
          32084 => x"80", -- $07d54
          32085 => x"7f", -- $07d55
          32086 => x"7f", -- $07d56
          32087 => x"7f", -- $07d57
          32088 => x"7f", -- $07d58
          32089 => x"7e", -- $07d59
          32090 => x"7e", -- $07d5a
          32091 => x"7e", -- $07d5b
          32092 => x"7e", -- $07d5c
          32093 => x"7e", -- $07d5d
          32094 => x"7e", -- $07d5e
          32095 => x"7e", -- $07d5f
          32096 => x"7e", -- $07d60
          32097 => x"7e", -- $07d61
          32098 => x"7e", -- $07d62
          32099 => x"7e", -- $07d63
          32100 => x"7f", -- $07d64
          32101 => x"7f", -- $07d65
          32102 => x"7f", -- $07d66
          32103 => x"7f", -- $07d67
          32104 => x"7f", -- $07d68
          32105 => x"7f", -- $07d69
          32106 => x"80", -- $07d6a
          32107 => x"80", -- $07d6b
          32108 => x"80", -- $07d6c
          32109 => x"80", -- $07d6d
          32110 => x"80", -- $07d6e
          32111 => x"80", -- $07d6f
          32112 => x"80", -- $07d70
          32113 => x"80", -- $07d71
          32114 => x"80", -- $07d72
          32115 => x"80", -- $07d73
          32116 => x"80", -- $07d74
          32117 => x"80", -- $07d75
          32118 => x"7f", -- $07d76
          32119 => x"7f", -- $07d77
          32120 => x"7f", -- $07d78
          32121 => x"7f", -- $07d79
          32122 => x"7f", -- $07d7a
          32123 => x"7f", -- $07d7b
          32124 => x"7f", -- $07d7c
          32125 => x"7f", -- $07d7d
          32126 => x"7f", -- $07d7e
          32127 => x"7f", -- $07d7f
          32128 => x"7f", -- $07d80
          32129 => x"7f", -- $07d81
          32130 => x"7f", -- $07d82
          32131 => x"7f", -- $07d83
          32132 => x"7f", -- $07d84
          32133 => x"7f", -- $07d85
          32134 => x"7f", -- $07d86
          32135 => x"7f", -- $07d87
          32136 => x"80", -- $07d88
          32137 => x"80", -- $07d89
          32138 => x"80", -- $07d8a
          32139 => x"80", -- $07d8b
          32140 => x"80", -- $07d8c
          32141 => x"80", -- $07d8d
          32142 => x"80", -- $07d8e
          32143 => x"80", -- $07d8f
          32144 => x"80", -- $07d90
          32145 => x"80", -- $07d91
          32146 => x"80", -- $07d92
          32147 => x"80", -- $07d93
          32148 => x"80", -- $07d94
          32149 => x"80", -- $07d95
          32150 => x"80", -- $07d96
          32151 => x"80", -- $07d97
          32152 => x"80", -- $07d98
          32153 => x"80", -- $07d99
          32154 => x"7f", -- $07d9a
          32155 => x"7f", -- $07d9b
          32156 => x"7f", -- $07d9c
          32157 => x"7f", -- $07d9d
          32158 => x"7f", -- $07d9e
          32159 => x"7f", -- $07d9f
          32160 => x"7f", -- $07da0
          32161 => x"7f", -- $07da1
          32162 => x"80", -- $07da2
          32163 => x"80", -- $07da3
          32164 => x"80", -- $07da4
          32165 => x"80", -- $07da5
          32166 => x"80", -- $07da6
          32167 => x"80", -- $07da7
          32168 => x"80", -- $07da8
          32169 => x"80", -- $07da9
          32170 => x"80", -- $07daa
          32171 => x"80", -- $07dab
          32172 => x"80", -- $07dac
          32173 => x"81", -- $07dad
          32174 => x"81", -- $07dae
          32175 => x"81", -- $07daf
          32176 => x"81", -- $07db0
          32177 => x"81", -- $07db1
          32178 => x"81", -- $07db2
          32179 => x"80", -- $07db3
          32180 => x"80", -- $07db4
          32181 => x"80", -- $07db5
          32182 => x"80", -- $07db6
          32183 => x"80", -- $07db7
          32184 => x"80", -- $07db8
          32185 => x"80", -- $07db9
          32186 => x"80", -- $07dba
          32187 => x"80", -- $07dbb
          32188 => x"80", -- $07dbc
          32189 => x"80", -- $07dbd
          32190 => x"80", -- $07dbe
          32191 => x"80", -- $07dbf
          32192 => x"80", -- $07dc0
          32193 => x"80", -- $07dc1
          32194 => x"80", -- $07dc2
          32195 => x"80", -- $07dc3
          32196 => x"80", -- $07dc4
          32197 => x"80", -- $07dc5
          32198 => x"80", -- $07dc6
          32199 => x"80", -- $07dc7
          32200 => x"80", -- $07dc8
          32201 => x"81", -- $07dc9
          32202 => x"81", -- $07dca
          32203 => x"81", -- $07dcb
          32204 => x"81", -- $07dcc
          32205 => x"82", -- $07dcd
          32206 => x"81", -- $07dce
          32207 => x"81", -- $07dcf
          32208 => x"81", -- $07dd0
          32209 => x"81", -- $07dd1
          32210 => x"81", -- $07dd2
          32211 => x"81", -- $07dd3
          32212 => x"81", -- $07dd4
          32213 => x"81", -- $07dd5
          32214 => x"81", -- $07dd6
          32215 => x"80", -- $07dd7
          32216 => x"80", -- $07dd8
          32217 => x"80", -- $07dd9
          32218 => x"80", -- $07dda
          32219 => x"80", -- $07ddb
          32220 => x"80", -- $07ddc
          32221 => x"80", -- $07ddd
          32222 => x"80", -- $07dde
          32223 => x"80", -- $07ddf
          32224 => x"80", -- $07de0
          32225 => x"80", -- $07de1
          32226 => x"80", -- $07de2
          32227 => x"80", -- $07de3
          32228 => x"80", -- $07de4
          32229 => x"81", -- $07de5
          32230 => x"81", -- $07de6
          32231 => x"81", -- $07de7
          32232 => x"81", -- $07de8
          32233 => x"82", -- $07de9
          32234 => x"82", -- $07dea
          32235 => x"81", -- $07deb
          32236 => x"82", -- $07dec
          32237 => x"82", -- $07ded
          32238 => x"82", -- $07dee
          32239 => x"82", -- $07def
          32240 => x"82", -- $07df0
          32241 => x"82", -- $07df1
          32242 => x"82", -- $07df2
          32243 => x"82", -- $07df3
          32244 => x"82", -- $07df4
          32245 => x"81", -- $07df5
          32246 => x"81", -- $07df6
          32247 => x"81", -- $07df7
          32248 => x"81", -- $07df8
          32249 => x"81", -- $07df9
          32250 => x"80", -- $07dfa
          32251 => x"80", -- $07dfb
          32252 => x"80", -- $07dfc
          32253 => x"80", -- $07dfd
          32254 => x"80", -- $07dfe
          32255 => x"80", -- $07dff
          32256 => x"80", -- $07e00
          32257 => x"80", -- $07e01
          32258 => x"80", -- $07e02
          32259 => x"81", -- $07e03
          32260 => x"81", -- $07e04
          32261 => x"81", -- $07e05
          32262 => x"81", -- $07e06
          32263 => x"82", -- $07e07
          32264 => x"82", -- $07e08
          32265 => x"82", -- $07e09
          32266 => x"82", -- $07e0a
          32267 => x"83", -- $07e0b
          32268 => x"83", -- $07e0c
          32269 => x"83", -- $07e0d
          32270 => x"83", -- $07e0e
          32271 => x"83", -- $07e0f
          32272 => x"83", -- $07e10
          32273 => x"83", -- $07e11
          32274 => x"83", -- $07e12
          32275 => x"82", -- $07e13
          32276 => x"82", -- $07e14
          32277 => x"82", -- $07e15
          32278 => x"82", -- $07e16
          32279 => x"81", -- $07e17
          32280 => x"81", -- $07e18
          32281 => x"81", -- $07e19
          32282 => x"81", -- $07e1a
          32283 => x"81", -- $07e1b
          32284 => x"81", -- $07e1c
          32285 => x"81", -- $07e1d
          32286 => x"81", -- $07e1e
          32287 => x"81", -- $07e1f
          32288 => x"81", -- $07e20
          32289 => x"81", -- $07e21
          32290 => x"81", -- $07e22
          32291 => x"81", -- $07e23
          32292 => x"81", -- $07e24
          32293 => x"81", -- $07e25
          32294 => x"82", -- $07e26
          32295 => x"82", -- $07e27
          32296 => x"82", -- $07e28
          32297 => x"82", -- $07e29
          32298 => x"83", -- $07e2a
          32299 => x"83", -- $07e2b
          32300 => x"83", -- $07e2c
          32301 => x"83", -- $07e2d
          32302 => x"83", -- $07e2e
          32303 => x"83", -- $07e2f
          32304 => x"83", -- $07e30
          32305 => x"83", -- $07e31
          32306 => x"83", -- $07e32
          32307 => x"83", -- $07e33
          32308 => x"83", -- $07e34
          32309 => x"82", -- $07e35
          32310 => x"82", -- $07e36
          32311 => x"82", -- $07e37
          32312 => x"81", -- $07e38
          32313 => x"81", -- $07e39
          32314 => x"81", -- $07e3a
          32315 => x"81", -- $07e3b
          32316 => x"80", -- $07e3c
          32317 => x"80", -- $07e3d
          32318 => x"80", -- $07e3e
          32319 => x"81", -- $07e3f
          32320 => x"81", -- $07e40
          32321 => x"81", -- $07e41
          32322 => x"81", -- $07e42
          32323 => x"81", -- $07e43
          32324 => x"81", -- $07e44
          32325 => x"81", -- $07e45
          32326 => x"81", -- $07e46
          32327 => x"82", -- $07e47
          32328 => x"82", -- $07e48
          32329 => x"82", -- $07e49
          32330 => x"82", -- $07e4a
          32331 => x"82", -- $07e4b
          32332 => x"83", -- $07e4c
          32333 => x"83", -- $07e4d
          32334 => x"83", -- $07e4e
          32335 => x"83", -- $07e4f
          32336 => x"83", -- $07e50
          32337 => x"83", -- $07e51
          32338 => x"82", -- $07e52
          32339 => x"82", -- $07e53
          32340 => x"82", -- $07e54
          32341 => x"81", -- $07e55
          32342 => x"81", -- $07e56
          32343 => x"81", -- $07e57
          32344 => x"81", -- $07e58
          32345 => x"81", -- $07e59
          32346 => x"80", -- $07e5a
          32347 => x"80", -- $07e5b
          32348 => x"80", -- $07e5c
          32349 => x"80", -- $07e5d
          32350 => x"80", -- $07e5e
          32351 => x"80", -- $07e5f
          32352 => x"80", -- $07e60
          32353 => x"80", -- $07e61
          32354 => x"80", -- $07e62
          32355 => x"80", -- $07e63
          32356 => x"81", -- $07e64
          32357 => x"81", -- $07e65
          32358 => x"81", -- $07e66
          32359 => x"82", -- $07e67
          32360 => x"82", -- $07e68
          32361 => x"82", -- $07e69
          32362 => x"82", -- $07e6a
          32363 => x"82", -- $07e6b
          32364 => x"83", -- $07e6c
          32365 => x"82", -- $07e6d
          32366 => x"83", -- $07e6e
          32367 => x"83", -- $07e6f
          32368 => x"82", -- $07e70
          32369 => x"82", -- $07e71
          32370 => x"82", -- $07e72
          32371 => x"82", -- $07e73
          32372 => x"82", -- $07e74
          32373 => x"82", -- $07e75
          32374 => x"81", -- $07e76
          32375 => x"81", -- $07e77
          32376 => x"81", -- $07e78
          32377 => x"81", -- $07e79
          32378 => x"80", -- $07e7a
          32379 => x"80", -- $07e7b
          32380 => x"80", -- $07e7c
          32381 => x"80", -- $07e7d
          32382 => x"80", -- $07e7e
          32383 => x"80", -- $07e7f
          32384 => x"80", -- $07e80
          32385 => x"80", -- $07e81
          32386 => x"81", -- $07e82
          32387 => x"81", -- $07e83
          32388 => x"81", -- $07e84
          32389 => x"81", -- $07e85
          32390 => x"82", -- $07e86
          32391 => x"82", -- $07e87
          32392 => x"82", -- $07e88
          32393 => x"82", -- $07e89
          32394 => x"82", -- $07e8a
          32395 => x"82", -- $07e8b
          32396 => x"83", -- $07e8c
          32397 => x"83", -- $07e8d
          32398 => x"83", -- $07e8e
          32399 => x"83", -- $07e8f
          32400 => x"83", -- $07e90
          32401 => x"82", -- $07e91
          32402 => x"82", -- $07e92
          32403 => x"82", -- $07e93
          32404 => x"82", -- $07e94
          32405 => x"82", -- $07e95
          32406 => x"81", -- $07e96
          32407 => x"81", -- $07e97
          32408 => x"81", -- $07e98
          32409 => x"81", -- $07e99
          32410 => x"81", -- $07e9a
          32411 => x"81", -- $07e9b
          32412 => x"81", -- $07e9c
          32413 => x"81", -- $07e9d
          32414 => x"81", -- $07e9e
          32415 => x"81", -- $07e9f
          32416 => x"81", -- $07ea0
          32417 => x"81", -- $07ea1
          32418 => x"81", -- $07ea2
          32419 => x"82", -- $07ea3
          32420 => x"82", -- $07ea4
          32421 => x"82", -- $07ea5
          32422 => x"82", -- $07ea6
          32423 => x"83", -- $07ea7
          32424 => x"83", -- $07ea8
          32425 => x"83", -- $07ea9
          32426 => x"83", -- $07eaa
          32427 => x"83", -- $07eab
          32428 => x"83", -- $07eac
          32429 => x"83", -- $07ead
          32430 => x"83", -- $07eae
          32431 => x"83", -- $07eaf
          32432 => x"83", -- $07eb0
          32433 => x"83", -- $07eb1
          32434 => x"83", -- $07eb2
          32435 => x"82", -- $07eb3
          32436 => x"82", -- $07eb4
          32437 => x"82", -- $07eb5
          32438 => x"82", -- $07eb6
          32439 => x"81", -- $07eb7
          32440 => x"81", -- $07eb8
          32441 => x"81", -- $07eb9
          32442 => x"81", -- $07eba
          32443 => x"81", -- $07ebb
          32444 => x"81", -- $07ebc
          32445 => x"81", -- $07ebd
          32446 => x"81", -- $07ebe
          32447 => x"81", -- $07ebf
          32448 => x"81", -- $07ec0
          32449 => x"82", -- $07ec1
          32450 => x"82", -- $07ec2
          32451 => x"82", -- $07ec3
          32452 => x"82", -- $07ec4
          32453 => x"83", -- $07ec5
          32454 => x"83", -- $07ec6
          32455 => x"83", -- $07ec7
          32456 => x"83", -- $07ec8
          32457 => x"83", -- $07ec9
          32458 => x"83", -- $07eca
          32459 => x"83", -- $07ecb
          32460 => x"83", -- $07ecc
          32461 => x"83", -- $07ecd
          32462 => x"83", -- $07ece
          32463 => x"83", -- $07ecf
          32464 => x"83", -- $07ed0
          32465 => x"83", -- $07ed1
          32466 => x"82", -- $07ed2
          32467 => x"82", -- $07ed3
          32468 => x"82", -- $07ed4
          32469 => x"82", -- $07ed5
          32470 => x"81", -- $07ed6
          32471 => x"81", -- $07ed7
          32472 => x"81", -- $07ed8
          32473 => x"81", -- $07ed9
          32474 => x"80", -- $07eda
          32475 => x"80", -- $07edb
          32476 => x"80", -- $07edc
          32477 => x"81", -- $07edd
          32478 => x"81", -- $07ede
          32479 => x"81", -- $07edf
          32480 => x"81", -- $07ee0
          32481 => x"81", -- $07ee1
          32482 => x"81", -- $07ee2
          32483 => x"81", -- $07ee3
          32484 => x"82", -- $07ee4
          32485 => x"82", -- $07ee5
          32486 => x"82", -- $07ee6
          32487 => x"82", -- $07ee7
          32488 => x"82", -- $07ee8
          32489 => x"82", -- $07ee9
          32490 => x"82", -- $07eea
          32491 => x"82", -- $07eeb
          32492 => x"82", -- $07eec
          32493 => x"82", -- $07eed
          32494 => x"82", -- $07eee
          32495 => x"81", -- $07eef
          32496 => x"81", -- $07ef0
          32497 => x"81", -- $07ef1
          32498 => x"81", -- $07ef2
          32499 => x"80", -- $07ef3
          32500 => x"80", -- $07ef4
          32501 => x"80", -- $07ef5
          32502 => x"80", -- $07ef6
          32503 => x"80", -- $07ef7
          32504 => x"80", -- $07ef8
          32505 => x"80", -- $07ef9
          32506 => x"80", -- $07efa
          32507 => x"80", -- $07efb
          32508 => x"80", -- $07efc
          32509 => x"80", -- $07efd
          32510 => x"80", -- $07efe
          32511 => x"80", -- $07eff
          32512 => x"80", -- $07f00
          32513 => x"80", -- $07f01
          32514 => x"80", -- $07f02
          32515 => x"80", -- $07f03
          32516 => x"81", -- $07f04
          32517 => x"81", -- $07f05
          32518 => x"81", -- $07f06
          32519 => x"81", -- $07f07
          32520 => x"81", -- $07f08
          32521 => x"81", -- $07f09
          32522 => x"80", -- $07f0a
          32523 => x"80", -- $07f0b
          32524 => x"80", -- $07f0c
          32525 => x"80", -- $07f0d
          32526 => x"80", -- $07f0e
          32527 => x"80", -- $07f0f
          32528 => x"80", -- $07f10
          32529 => x"80", -- $07f11
          32530 => x"80", -- $07f12
          32531 => x"80", -- $07f13
          32532 => x"80", -- $07f14
          32533 => x"80", -- $07f15
          32534 => x"7f", -- $07f16
          32535 => x"7f", -- $07f17
          32536 => x"7f", -- $07f18
          32537 => x"7f", -- $07f19
          32538 => x"7f", -- $07f1a
          32539 => x"7f", -- $07f1b
          32540 => x"7f", -- $07f1c
          32541 => x"7f", -- $07f1d
          32542 => x"80", -- $07f1e
          32543 => x"80", -- $07f1f
          32544 => x"80", -- $07f20
          32545 => x"80", -- $07f21
          32546 => x"80", -- $07f22
          32547 => x"80", -- $07f23
          32548 => x"80", -- $07f24
          32549 => x"80", -- $07f25
          32550 => x"80", -- $07f26
          32551 => x"80", -- $07f27
          32552 => x"80", -- $07f28
          32553 => x"80", -- $07f29
          32554 => x"80", -- $07f2a
          32555 => x"80", -- $07f2b
          32556 => x"80", -- $07f2c
          32557 => x"80", -- $07f2d
          32558 => x"80", -- $07f2e
          32559 => x"80", -- $07f2f
          32560 => x"7f", -- $07f30
          32561 => x"7f", -- $07f31
          32562 => x"7f", -- $07f32
          32563 => x"7f", -- $07f33
          32564 => x"7f", -- $07f34
          32565 => x"7f", -- $07f35
          32566 => x"7f", -- $07f36
          32567 => x"7e", -- $07f37
          32568 => x"7e", -- $07f38
          32569 => x"7f", -- $07f39
          32570 => x"7f", -- $07f3a
          32571 => x"7f", -- $07f3b
          32572 => x"7f", -- $07f3c
          32573 => x"7f", -- $07f3d
          32574 => x"7f", -- $07f3e
          32575 => x"7f", -- $07f3f
          32576 => x"7f", -- $07f40
          32577 => x"80", -- $07f41
          32578 => x"80", -- $07f42
          32579 => x"80", -- $07f43
          32580 => x"80", -- $07f44
          32581 => x"80", -- $07f45
          32582 => x"80", -- $07f46
          32583 => x"80", -- $07f47
          32584 => x"80", -- $07f48
          32585 => x"80", -- $07f49
          32586 => x"80", -- $07f4a
          32587 => x"80", -- $07f4b
          32588 => x"7f", -- $07f4c
          32589 => x"7f", -- $07f4d
          32590 => x"7f", -- $07f4e
          32591 => x"7f", -- $07f4f
          32592 => x"7f", -- $07f50
          32593 => x"7f", -- $07f51
          32594 => x"7f", -- $07f52
          32595 => x"7f", -- $07f53
          32596 => x"7f", -- $07f54
          32597 => x"7f", -- $07f55
          32598 => x"7f", -- $07f56
          32599 => x"7f", -- $07f57
          32600 => x"7f", -- $07f58
          32601 => x"7f", -- $07f59
          32602 => x"7f", -- $07f5a
          32603 => x"7f", -- $07f5b
          32604 => x"7f", -- $07f5c
          32605 => x"7f", -- $07f5d
          32606 => x"7f", -- $07f5e
          32607 => x"80", -- $07f5f
          32608 => x"80", -- $07f60
          32609 => x"80", -- $07f61
          32610 => x"80", -- $07f62
          32611 => x"80", -- $07f63
          32612 => x"80", -- $07f64
          32613 => x"80", -- $07f65
          32614 => x"80", -- $07f66
          32615 => x"80", -- $07f67
          32616 => x"80", -- $07f68
          32617 => x"80", -- $07f69
          32618 => x"7f", -- $07f6a
          32619 => x"7f", -- $07f6b
          32620 => x"7f", -- $07f6c
          32621 => x"7f", -- $07f6d
          32622 => x"7f", -- $07f6e
          32623 => x"7f", -- $07f6f
          32624 => x"7f", -- $07f70
          32625 => x"7f", -- $07f71
          32626 => x"7f", -- $07f72
          32627 => x"7f", -- $07f73
          32628 => x"7e", -- $07f74
          32629 => x"7e", -- $07f75
          32630 => x"7f", -- $07f76
          32631 => x"7f", -- $07f77
          32632 => x"7f", -- $07f78
          32633 => x"7f", -- $07f79
          32634 => x"7f", -- $07f7a
          32635 => x"7f", -- $07f7b
          32636 => x"80", -- $07f7c
          32637 => x"80", -- $07f7d
          32638 => x"80", -- $07f7e
          32639 => x"80", -- $07f7f
          32640 => x"80", -- $07f80
          32641 => x"80", -- $07f81
          32642 => x"80", -- $07f82
          32643 => x"80", -- $07f83
          32644 => x"80", -- $07f84
          32645 => x"80", -- $07f85
          32646 => x"80", -- $07f86
          32647 => x"80", -- $07f87
          32648 => x"80", -- $07f88
          32649 => x"7f", -- $07f89
          32650 => x"7f", -- $07f8a
          32651 => x"7f", -- $07f8b
          32652 => x"7f", -- $07f8c
          32653 => x"7f", -- $07f8d
          32654 => x"7f", -- $07f8e
          32655 => x"7f", -- $07f8f
          32656 => x"7e", -- $07f90
          32657 => x"7f", -- $07f91
          32658 => x"7e", -- $07f92
          32659 => x"7e", -- $07f93
          32660 => x"7f", -- $07f94
          32661 => x"7f", -- $07f95
          32662 => x"7f", -- $07f96
          32663 => x"7f", -- $07f97
          32664 => x"7f", -- $07f98
          32665 => x"7f", -- $07f99
          32666 => x"7f", -- $07f9a
          32667 => x"7f", -- $07f9b
          32668 => x"7f", -- $07f9c
          32669 => x"7f", -- $07f9d
          32670 => x"7f", -- $07f9e
          32671 => x"80", -- $07f9f
          32672 => x"80", -- $07fa0
          32673 => x"80", -- $07fa1
          32674 => x"80", -- $07fa2
          32675 => x"7f", -- $07fa3
          32676 => x"7f", -- $07fa4
          32677 => x"7f", -- $07fa5
          32678 => x"7f", -- $07fa6
          32679 => x"7f", -- $07fa7
          32680 => x"7f", -- $07fa8
          32681 => x"7f", -- $07fa9
          32682 => x"7f", -- $07faa
          32683 => x"7e", -- $07fab
          32684 => x"7e", -- $07fac
          32685 => x"7e", -- $07fad
          32686 => x"7e", -- $07fae
          32687 => x"7e", -- $07faf
          32688 => x"7e", -- $07fb0
          32689 => x"7e", -- $07fb1
          32690 => x"7e", -- $07fb2
          32691 => x"7e", -- $07fb3
          32692 => x"7e", -- $07fb4
          32693 => x"7e", -- $07fb5
          32694 => x"7e", -- $07fb6
          32695 => x"7f", -- $07fb7
          32696 => x"7f", -- $07fb8
          32697 => x"7f", -- $07fb9
          32698 => x"7f", -- $07fba
          32699 => x"7f", -- $07fbb
          32700 => x"7f", -- $07fbc
          32701 => x"7f", -- $07fbd
          32702 => x"7f", -- $07fbe
          32703 => x"7f", -- $07fbf
          32704 => x"7f", -- $07fc0
          32705 => x"7f", -- $07fc1
          32706 => x"7f", -- $07fc2
          32707 => x"7f", -- $07fc3
          32708 => x"7f", -- $07fc4
          32709 => x"7f", -- $07fc5
          32710 => x"7f", -- $07fc6
          32711 => x"7e", -- $07fc7
          32712 => x"7e", -- $07fc8
          32713 => x"7e", -- $07fc9
          32714 => x"7e", -- $07fca
          32715 => x"7e", -- $07fcb
          32716 => x"7e", -- $07fcc
          32717 => x"7e", -- $07fcd
          32718 => x"7e", -- $07fce
          32719 => x"7e", -- $07fcf
          32720 => x"7e", -- $07fd0
          32721 => x"7e", -- $07fd1
          32722 => x"7e", -- $07fd2
          32723 => x"7e", -- $07fd3
          32724 => x"7e", -- $07fd4
          32725 => x"7e", -- $07fd5
          32726 => x"7e", -- $07fd6
          32727 => x"7e", -- $07fd7
          32728 => x"7e", -- $07fd8
          32729 => x"7f", -- $07fd9
          32730 => x"7f", -- $07fda
          32731 => x"7f", -- $07fdb
          32732 => x"7f", -- $07fdc
          32733 => x"7f", -- $07fdd
          32734 => x"7f", -- $07fde
          32735 => x"7f", -- $07fdf
          32736 => x"7f", -- $07fe0
          32737 => x"7f", -- $07fe1
          32738 => x"7f", -- $07fe2
          32739 => x"7f", -- $07fe3
          32740 => x"7e", -- $07fe4
          32741 => x"7e", -- $07fe5
          32742 => x"7e", -- $07fe6
          32743 => x"7e", -- $07fe7
          32744 => x"7e", -- $07fe8
          32745 => x"7e", -- $07fe9
          32746 => x"7d", -- $07fea
          32747 => x"7d", -- $07feb
          32748 => x"7d", -- $07fec
          32749 => x"7d", -- $07fed
          32750 => x"7d", -- $07fee
          32751 => x"7d", -- $07fef
          32752 => x"7d", -- $07ff0
          32753 => x"7d", -- $07ff1
          32754 => x"7e", -- $07ff2
          32755 => x"7e", -- $07ff3
          32756 => x"7e", -- $07ff4
          32757 => x"7e", -- $07ff5
          32758 => x"7e", -- $07ff6
          32759 => x"7e", -- $07ff7
          32760 => x"7e", -- $07ff8
          32761 => x"7e", -- $07ff9
          32762 => x"7e", -- $07ffa
          32763 => x"7e", -- $07ffb
          32764 => x"7f", -- $07ffc
          32765 => x"7f", -- $07ffd
          32766 => x"7f", -- $07ffe
          32767 => x"7f", -- $07fff
          32768 => x"7e", -- $08000
          32769 => x"7e", -- $08001
          32770 => x"7e", -- $08002
          32771 => x"7e", -- $08003
          32772 => x"7e", -- $08004
          32773 => x"7e", -- $08005
          32774 => x"7e", -- $08006
          32775 => x"7d", -- $08007
          32776 => x"7d", -- $08008
          32777 => x"7d", -- $08009
          32778 => x"7d", -- $0800a
          32779 => x"7d", -- $0800b
          32780 => x"7d", -- $0800c
          32781 => x"7d", -- $0800d
          32782 => x"7d", -- $0800e
          32783 => x"7d", -- $0800f
          32784 => x"7d", -- $08010
          32785 => x"7e", -- $08011
          32786 => x"7e", -- $08012
          32787 => x"7e", -- $08013
          32788 => x"7e", -- $08014
          32789 => x"7e", -- $08015
          32790 => x"7e", -- $08016
          32791 => x"7f", -- $08017
          32792 => x"7f", -- $08018
          32793 => x"7f", -- $08019
          32794 => x"7f", -- $0801a
          32795 => x"7f", -- $0801b
          32796 => x"7f", -- $0801c
          32797 => x"7f", -- $0801d
          32798 => x"7f", -- $0801e
          32799 => x"7f", -- $0801f
          32800 => x"7f", -- $08020
          32801 => x"7e", -- $08021
          32802 => x"7e", -- $08022
          32803 => x"7e", -- $08023
          32804 => x"7e", -- $08024
          32805 => x"7e", -- $08025
          32806 => x"7e", -- $08026
          32807 => x"7e", -- $08027
          32808 => x"7e", -- $08028
          32809 => x"7e", -- $08029
          32810 => x"7e", -- $0802a
          32811 => x"7e", -- $0802b
          32812 => x"7d", -- $0802c
          32813 => x"7e", -- $0802d
          32814 => x"7e", -- $0802e
          32815 => x"7e", -- $0802f
          32816 => x"7e", -- $08030
          32817 => x"7e", -- $08031
          32818 => x"7e", -- $08032
          32819 => x"7f", -- $08033
          32820 => x"7f", -- $08034
          32821 => x"7f", -- $08035
          32822 => x"7f", -- $08036
          32823 => x"7f", -- $08037
          32824 => x"7f", -- $08038
          32825 => x"7f", -- $08039
          32826 => x"7f", -- $0803a
          32827 => x"7f", -- $0803b
          32828 => x"7f", -- $0803c
          32829 => x"7f", -- $0803d
          32830 => x"7f", -- $0803e
          32831 => x"7f", -- $0803f
          32832 => x"7f", -- $08040
          32833 => x"7f", -- $08041
          32834 => x"7f", -- $08042
          32835 => x"7f", -- $08043
          32836 => x"7e", -- $08044
          32837 => x"7e", -- $08045
          32838 => x"7e", -- $08046
          32839 => x"7e", -- $08047
          32840 => x"7e", -- $08048
          32841 => x"7e", -- $08049
          32842 => x"7e", -- $0804a
          32843 => x"7e", -- $0804b
          32844 => x"7e", -- $0804c
          32845 => x"7e", -- $0804d
          32846 => x"7e", -- $0804e
          32847 => x"7f", -- $0804f
          32848 => x"7f", -- $08050
          32849 => x"7f", -- $08051
          32850 => x"7f", -- $08052
          32851 => x"7f", -- $08053
          32852 => x"7f", -- $08054
          32853 => x"80", -- $08055
          32854 => x"80", -- $08056
          32855 => x"80", -- $08057
          32856 => x"80", -- $08058
          32857 => x"80", -- $08059
          32858 => x"80", -- $0805a
          32859 => x"80", -- $0805b
          32860 => x"80", -- $0805c
          32861 => x"80", -- $0805d
          32862 => x"80", -- $0805e
          32863 => x"80", -- $0805f
          32864 => x"7f", -- $08060
          32865 => x"7f", -- $08061
          32866 => x"7f", -- $08062
          32867 => x"7f", -- $08063
          32868 => x"7f", -- $08064
          32869 => x"7f", -- $08065
          32870 => x"7f", -- $08066
          32871 => x"7f", -- $08067
          32872 => x"7f", -- $08068
          32873 => x"7f", -- $08069
          32874 => x"7f", -- $0806a
          32875 => x"7f", -- $0806b
          32876 => x"7f", -- $0806c
          32877 => x"7f", -- $0806d
          32878 => x"7f", -- $0806e
          32879 => x"7f", -- $0806f
          32880 => x"80", -- $08070
          32881 => x"80", -- $08071
          32882 => x"80", -- $08072
          32883 => x"80", -- $08073
          32884 => x"80", -- $08074
          32885 => x"80", -- $08075
          32886 => x"80", -- $08076
          32887 => x"80", -- $08077
          32888 => x"80", -- $08078
          32889 => x"80", -- $08079
          32890 => x"80", -- $0807a
          32891 => x"80", -- $0807b
          32892 => x"80", -- $0807c
          32893 => x"80", -- $0807d
          32894 => x"80", -- $0807e
          32895 => x"80", -- $0807f
          32896 => x"80", -- $08080
          32897 => x"80", -- $08081
          32898 => x"80", -- $08082
          32899 => x"80", -- $08083
          32900 => x"80", -- $08084
          32901 => x"80", -- $08085
          32902 => x"80", -- $08086
          32903 => x"80", -- $08087
          32904 => x"80", -- $08088
          32905 => x"80", -- $08089
          32906 => x"80", -- $0808a
          32907 => x"80", -- $0808b
          32908 => x"80", -- $0808c
          32909 => x"80", -- $0808d
          32910 => x"80", -- $0808e
          32911 => x"80", -- $0808f
          32912 => x"80", -- $08090
          32913 => x"80", -- $08091
          32914 => x"80", -- $08092
          32915 => x"80", -- $08093
          32916 => x"81", -- $08094
          32917 => x"81", -- $08095
          32918 => x"81", -- $08096
          32919 => x"81", -- $08097
          32920 => x"81", -- $08098
          32921 => x"81", -- $08099
          32922 => x"81", -- $0809a
          32923 => x"81", -- $0809b
          32924 => x"80", -- $0809c
          32925 => x"80", -- $0809d
          32926 => x"80", -- $0809e
          32927 => x"80", -- $0809f
          32928 => x"80", -- $080a0
          32929 => x"80", -- $080a1
          32930 => x"80", -- $080a2
          32931 => x"80", -- $080a3
          32932 => x"80", -- $080a4
          32933 => x"80", -- $080a5
          32934 => x"80", -- $080a6
          32935 => x"80", -- $080a7
          32936 => x"80", -- $080a8
          32937 => x"80", -- $080a9
          32938 => x"80", -- $080aa
          32939 => x"80", -- $080ab
          32940 => x"80", -- $080ac
          32941 => x"80", -- $080ad
          32942 => x"80", -- $080ae
          32943 => x"80", -- $080af
          32944 => x"80", -- $080b0
          32945 => x"81", -- $080b1
          32946 => x"81", -- $080b2
          32947 => x"81", -- $080b3
          32948 => x"81", -- $080b4
          32949 => x"81", -- $080b5
          32950 => x"81", -- $080b6
          32951 => x"81", -- $080b7
          32952 => x"81", -- $080b8
          32953 => x"81", -- $080b9
          32954 => x"81", -- $080ba
          32955 => x"80", -- $080bb
          32956 => x"80", -- $080bc
          32957 => x"80", -- $080bd
          32958 => x"80", -- $080be
          32959 => x"80", -- $080bf
          32960 => x"80", -- $080c0
          32961 => x"80", -- $080c1
          32962 => x"80", -- $080c2
          32963 => x"80", -- $080c3
          32964 => x"80", -- $080c4
          32965 => x"80", -- $080c5
          32966 => x"80", -- $080c6
          32967 => x"80", -- $080c7
          32968 => x"80", -- $080c8
          32969 => x"80", -- $080c9
          32970 => x"80", -- $080ca
          32971 => x"80", -- $080cb
          32972 => x"80", -- $080cc
          32973 => x"80", -- $080cd
          32974 => x"80", -- $080ce
          32975 => x"81", -- $080cf
          32976 => x"81", -- $080d0
          32977 => x"81", -- $080d1
          32978 => x"81", -- $080d2
          32979 => x"81", -- $080d3
          32980 => x"81", -- $080d4
          32981 => x"81", -- $080d5
          32982 => x"81", -- $080d6
          32983 => x"81", -- $080d7
          32984 => x"81", -- $080d8
          32985 => x"81", -- $080d9
          32986 => x"81", -- $080da
          32987 => x"81", -- $080db
          32988 => x"81", -- $080dc
          32989 => x"80", -- $080dd
          32990 => x"80", -- $080de
          32991 => x"80", -- $080df
          32992 => x"80", -- $080e0
          32993 => x"80", -- $080e1
          32994 => x"80", -- $080e2
          32995 => x"80", -- $080e3
          32996 => x"80", -- $080e4
          32997 => x"80", -- $080e5
          32998 => x"80", -- $080e6
          32999 => x"80", -- $080e7
          33000 => x"80", -- $080e8
          33001 => x"80", -- $080e9
          33002 => x"80", -- $080ea
          33003 => x"80", -- $080eb
          33004 => x"80", -- $080ec
          33005 => x"81", -- $080ed
          33006 => x"81", -- $080ee
          33007 => x"81", -- $080ef
          33008 => x"81", -- $080f0
          33009 => x"81", -- $080f1
          33010 => x"82", -- $080f2
          33011 => x"82", -- $080f3
          33012 => x"82", -- $080f4
          33013 => x"82", -- $080f5
          33014 => x"82", -- $080f6
          33015 => x"82", -- $080f7
          33016 => x"81", -- $080f8
          33017 => x"81", -- $080f9
          33018 => x"81", -- $080fa
          33019 => x"81", -- $080fb
          33020 => x"81", -- $080fc
          33021 => x"81", -- $080fd
          33022 => x"80", -- $080fe
          33023 => x"80", -- $080ff
          33024 => x"80", -- $08100
          33025 => x"80", -- $08101
          33026 => x"80", -- $08102
          33027 => x"80", -- $08103
          33028 => x"80", -- $08104
          33029 => x"80", -- $08105
          33030 => x"80", -- $08106
          33031 => x"80", -- $08107
          33032 => x"80", -- $08108
          33033 => x"81", -- $08109
          33034 => x"81", -- $0810a
          33035 => x"81", -- $0810b
          33036 => x"82", -- $0810c
          33037 => x"82", -- $0810d
          33038 => x"82", -- $0810e
          33039 => x"82", -- $0810f
          33040 => x"82", -- $08110
          33041 => x"83", -- $08111
          33042 => x"83", -- $08112
          33043 => x"83", -- $08113
          33044 => x"83", -- $08114
          33045 => x"83", -- $08115
          33046 => x"82", -- $08116
          33047 => x"82", -- $08117
          33048 => x"82", -- $08118
          33049 => x"82", -- $08119
          33050 => x"82", -- $0811a
          33051 => x"82", -- $0811b
          33052 => x"82", -- $0811c
          33053 => x"81", -- $0811d
          33054 => x"81", -- $0811e
          33055 => x"81", -- $0811f
          33056 => x"81", -- $08120
          33057 => x"81", -- $08121
          33058 => x"81", -- $08122
          33059 => x"81", -- $08123
          33060 => x"81", -- $08124
          33061 => x"81", -- $08125
          33062 => x"82", -- $08126
          33063 => x"82", -- $08127
          33064 => x"82", -- $08128
          33065 => x"82", -- $08129
          33066 => x"83", -- $0812a
          33067 => x"83", -- $0812b
          33068 => x"83", -- $0812c
          33069 => x"83", -- $0812d
          33070 => x"83", -- $0812e
          33071 => x"83", -- $0812f
          33072 => x"84", -- $08130
          33073 => x"83", -- $08131
          33074 => x"83", -- $08132
          33075 => x"84", -- $08133
          33076 => x"83", -- $08134
          33077 => x"83", -- $08135
          33078 => x"83", -- $08136
          33079 => x"83", -- $08137
          33080 => x"83", -- $08138
          33081 => x"83", -- $08139
          33082 => x"83", -- $0813a
          33083 => x"82", -- $0813b
          33084 => x"82", -- $0813c
          33085 => x"82", -- $0813d
          33086 => x"82", -- $0813e
          33087 => x"82", -- $0813f
          33088 => x"81", -- $08140
          33089 => x"82", -- $08141
          33090 => x"81", -- $08142
          33091 => x"82", -- $08143
          33092 => x"82", -- $08144
          33093 => x"82", -- $08145
          33094 => x"82", -- $08146
          33095 => x"82", -- $08147
          33096 => x"83", -- $08148
          33097 => x"83", -- $08149
          33098 => x"83", -- $0814a
          33099 => x"83", -- $0814b
          33100 => x"83", -- $0814c
          33101 => x"84", -- $0814d
          33102 => x"84", -- $0814e
          33103 => x"84", -- $0814f
          33104 => x"84", -- $08150
          33105 => x"84", -- $08151
          33106 => x"84", -- $08152
          33107 => x"84", -- $08153
          33108 => x"84", -- $08154
          33109 => x"84", -- $08155
          33110 => x"83", -- $08156
          33111 => x"83", -- $08157
          33112 => x"83", -- $08158
          33113 => x"83", -- $08159
          33114 => x"82", -- $0815a
          33115 => x"82", -- $0815b
          33116 => x"82", -- $0815c
          33117 => x"82", -- $0815d
          33118 => x"82", -- $0815e
          33119 => x"82", -- $0815f
          33120 => x"82", -- $08160
          33121 => x"81", -- $08161
          33122 => x"81", -- $08162
          33123 => x"81", -- $08163
          33124 => x"81", -- $08164
          33125 => x"81", -- $08165
          33126 => x"82", -- $08166
          33127 => x"82", -- $08167
          33128 => x"82", -- $08168
          33129 => x"83", -- $08169
          33130 => x"83", -- $0816a
          33131 => x"83", -- $0816b
          33132 => x"83", -- $0816c
          33133 => x"83", -- $0816d
          33134 => x"83", -- $0816e
          33135 => x"83", -- $0816f
          33136 => x"83", -- $08170
          33137 => x"83", -- $08171
          33138 => x"83", -- $08172
          33139 => x"83", -- $08173
          33140 => x"83", -- $08174
          33141 => x"83", -- $08175
          33142 => x"83", -- $08176
          33143 => x"82", -- $08177
          33144 => x"82", -- $08178
          33145 => x"82", -- $08179
          33146 => x"82", -- $0817a
          33147 => x"81", -- $0817b
          33148 => x"81", -- $0817c
          33149 => x"81", -- $0817d
          33150 => x"81", -- $0817e
          33151 => x"81", -- $0817f
          33152 => x"81", -- $08180
          33153 => x"81", -- $08181
          33154 => x"81", -- $08182
          33155 => x"81", -- $08183
          33156 => x"81", -- $08184
          33157 => x"81", -- $08185
          33158 => x"81", -- $08186
          33159 => x"81", -- $08187
          33160 => x"82", -- $08188
          33161 => x"82", -- $08189
          33162 => x"82", -- $0818a
          33163 => x"82", -- $0818b
          33164 => x"82", -- $0818c
          33165 => x"83", -- $0818d
          33166 => x"83", -- $0818e
          33167 => x"83", -- $0818f
          33168 => x"83", -- $08190
          33169 => x"83", -- $08191
          33170 => x"83", -- $08192
          33171 => x"83", -- $08193
          33172 => x"82", -- $08194
          33173 => x"82", -- $08195
          33174 => x"82", -- $08196
          33175 => x"82", -- $08197
          33176 => x"81", -- $08198
          33177 => x"81", -- $08199
          33178 => x"81", -- $0819a
          33179 => x"81", -- $0819b
          33180 => x"80", -- $0819c
          33181 => x"80", -- $0819d
          33182 => x"80", -- $0819e
          33183 => x"80", -- $0819f
          33184 => x"80", -- $081a0
          33185 => x"80", -- $081a1
          33186 => x"80", -- $081a2
          33187 => x"80", -- $081a3
          33188 => x"80", -- $081a4
          33189 => x"81", -- $081a5
          33190 => x"81", -- $081a6
          33191 => x"81", -- $081a7
          33192 => x"81", -- $081a8
          33193 => x"81", -- $081a9
          33194 => x"82", -- $081aa
          33195 => x"82", -- $081ab
          33196 => x"82", -- $081ac
          33197 => x"82", -- $081ad
          33198 => x"82", -- $081ae
          33199 => x"83", -- $081af
          33200 => x"83", -- $081b0
          33201 => x"82", -- $081b1
          33202 => x"82", -- $081b2
          33203 => x"82", -- $081b3
          33204 => x"82", -- $081b4
          33205 => x"82", -- $081b5
          33206 => x"82", -- $081b6
          33207 => x"81", -- $081b7
          33208 => x"81", -- $081b8
          33209 => x"81", -- $081b9
          33210 => x"81", -- $081ba
          33211 => x"80", -- $081bb
          33212 => x"80", -- $081bc
          33213 => x"80", -- $081bd
          33214 => x"80", -- $081be
          33215 => x"80", -- $081bf
          33216 => x"80", -- $081c0
          33217 => x"80", -- $081c1
          33218 => x"80", -- $081c2
          33219 => x"80", -- $081c3
          33220 => x"80", -- $081c4
          33221 => x"80", -- $081c5
          33222 => x"80", -- $081c6
          33223 => x"80", -- $081c7
          33224 => x"81", -- $081c8
          33225 => x"81", -- $081c9
          33226 => x"81", -- $081ca
          33227 => x"81", -- $081cb
          33228 => x"81", -- $081cc
          33229 => x"81", -- $081cd
          33230 => x"82", -- $081ce
          33231 => x"82", -- $081cf
          33232 => x"82", -- $081d0
          33233 => x"82", -- $081d1
          33234 => x"82", -- $081d2
          33235 => x"82", -- $081d3
          33236 => x"81", -- $081d4
          33237 => x"81", -- $081d5
          33238 => x"81", -- $081d6
          33239 => x"81", -- $081d7
          33240 => x"80", -- $081d8
          33241 => x"80", -- $081d9
          33242 => x"80", -- $081da
          33243 => x"80", -- $081db
          33244 => x"80", -- $081dc
          33245 => x"80", -- $081dd
          33246 => x"80", -- $081de
          33247 => x"80", -- $081df
          33248 => x"80", -- $081e0
          33249 => x"80", -- $081e1
          33250 => x"80", -- $081e2
          33251 => x"80", -- $081e3
          33252 => x"80", -- $081e4
          33253 => x"80", -- $081e5
          33254 => x"80", -- $081e6
          33255 => x"80", -- $081e7
          33256 => x"80", -- $081e8
          33257 => x"80", -- $081e9
          33258 => x"81", -- $081ea
          33259 => x"81", -- $081eb
          33260 => x"81", -- $081ec
          33261 => x"81", -- $081ed
          33262 => x"82", -- $081ee
          33263 => x"82", -- $081ef
          33264 => x"82", -- $081f0
          33265 => x"82", -- $081f1
          33266 => x"81", -- $081f2
          33267 => x"81", -- $081f3
          33268 => x"81", -- $081f4
          33269 => x"81", -- $081f5
          33270 => x"81", -- $081f6
          33271 => x"81", -- $081f7
          33272 => x"80", -- $081f8
          33273 => x"80", -- $081f9
          33274 => x"80", -- $081fa
          33275 => x"80", -- $081fb
          33276 => x"80", -- $081fc
          33277 => x"80", -- $081fd
          33278 => x"80", -- $081fe
          33279 => x"80", -- $081ff
          33280 => x"80", -- $08200
          33281 => x"80", -- $08201
          33282 => x"80", -- $08202
          33283 => x"80", -- $08203
          33284 => x"80", -- $08204
          33285 => x"80", -- $08205
          33286 => x"80", -- $08206
          33287 => x"80", -- $08207
          33288 => x"80", -- $08208
          33289 => x"80", -- $08209
          33290 => x"80", -- $0820a
          33291 => x"81", -- $0820b
          33292 => x"81", -- $0820c
          33293 => x"81", -- $0820d
          33294 => x"81", -- $0820e
          33295 => x"81", -- $0820f
          33296 => x"81", -- $08210
          33297 => x"81", -- $08211
          33298 => x"81", -- $08212
          33299 => x"81", -- $08213
          33300 => x"81", -- $08214
          33301 => x"81", -- $08215
          33302 => x"81", -- $08216
          33303 => x"81", -- $08217
          33304 => x"80", -- $08218
          33305 => x"80", -- $08219
          33306 => x"80", -- $0821a
          33307 => x"80", -- $0821b
          33308 => x"80", -- $0821c
          33309 => x"80", -- $0821d
          33310 => x"80", -- $0821e
          33311 => x"80", -- $0821f
          33312 => x"80", -- $08220
          33313 => x"80", -- $08221
          33314 => x"80", -- $08222
          33315 => x"80", -- $08223
          33316 => x"80", -- $08224
          33317 => x"80", -- $08225
          33318 => x"80", -- $08226
          33319 => x"80", -- $08227
          33320 => x"80", -- $08228
          33321 => x"80", -- $08229
          33322 => x"80", -- $0822a
          33323 => x"80", -- $0822b
          33324 => x"80", -- $0822c
          33325 => x"80", -- $0822d
          33326 => x"80", -- $0822e
          33327 => x"80", -- $0822f
          33328 => x"80", -- $08230
          33329 => x"80", -- $08231
          33330 => x"80", -- $08232
          33331 => x"80", -- $08233
          33332 => x"80", -- $08234
          33333 => x"80", -- $08235
          33334 => x"80", -- $08236
          33335 => x"80", -- $08237
          33336 => x"80", -- $08238
          33337 => x"80", -- $08239
          33338 => x"80", -- $0823a
          33339 => x"80", -- $0823b
          33340 => x"80", -- $0823c
          33341 => x"80", -- $0823d
          33342 => x"80", -- $0823e
          33343 => x"7f", -- $0823f
          33344 => x"7f", -- $08240
          33345 => x"7f", -- $08241
          33346 => x"7f", -- $08242
          33347 => x"7f", -- $08243
          33348 => x"7f", -- $08244
          33349 => x"7f", -- $08245
          33350 => x"7f", -- $08246
          33351 => x"7f", -- $08247
          33352 => x"7f", -- $08248
          33353 => x"80", -- $08249
          33354 => x"80", -- $0824a
          33355 => x"80", -- $0824b
          33356 => x"80", -- $0824c
          33357 => x"80", -- $0824d
          33358 => x"80", -- $0824e
          33359 => x"80", -- $0824f
          33360 => x"80", -- $08250
          33361 => x"80", -- $08251
          33362 => x"80", -- $08252
          33363 => x"80", -- $08253
          33364 => x"80", -- $08254
          33365 => x"80", -- $08255
          33366 => x"80", -- $08256
          33367 => x"80", -- $08257
          33368 => x"80", -- $08258
          33369 => x"80", -- $08259
          33370 => x"80", -- $0825a
          33371 => x"7f", -- $0825b
          33372 => x"7f", -- $0825c
          33373 => x"7f", -- $0825d
          33374 => x"7f", -- $0825e
          33375 => x"7f", -- $0825f
          33376 => x"7f", -- $08260
          33377 => x"7f", -- $08261
          33378 => x"7f", -- $08262
          33379 => x"7f", -- $08263
          33380 => x"7f", -- $08264
          33381 => x"7f", -- $08265
          33382 => x"7f", -- $08266
          33383 => x"7f", -- $08267
          33384 => x"7f", -- $08268
          33385 => x"7f", -- $08269
          33386 => x"7f", -- $0826a
          33387 => x"7f", -- $0826b
          33388 => x"7f", -- $0826c
          33389 => x"7f", -- $0826d
          33390 => x"7f", -- $0826e
          33391 => x"7f", -- $0826f
          33392 => x"7f", -- $08270
          33393 => x"7f", -- $08271
          33394 => x"7f", -- $08272
          33395 => x"7f", -- $08273
          33396 => x"7f", -- $08274
          33397 => x"7f", -- $08275
          33398 => x"7f", -- $08276
          33399 => x"7f", -- $08277
          33400 => x"7f", -- $08278
          33401 => x"7f", -- $08279
          33402 => x"7f", -- $0827a
          33403 => x"7f", -- $0827b
          33404 => x"7f", -- $0827c
          33405 => x"7f", -- $0827d
          33406 => x"7f", -- $0827e
          33407 => x"7f", -- $0827f
          33408 => x"7e", -- $08280
          33409 => x"7e", -- $08281
          33410 => x"7e", -- $08282
          33411 => x"7e", -- $08283
          33412 => x"7e", -- $08284
          33413 => x"7e", -- $08285
          33414 => x"7e", -- $08286
          33415 => x"7e", -- $08287
          33416 => x"7e", -- $08288
          33417 => x"7e", -- $08289
          33418 => x"7e", -- $0828a
          33419 => x"7e", -- $0828b
          33420 => x"7e", -- $0828c
          33421 => x"7e", -- $0828d
          33422 => x"7e", -- $0828e
          33423 => x"7e", -- $0828f
          33424 => x"7e", -- $08290
          33425 => x"7e", -- $08291
          33426 => x"7e", -- $08292
          33427 => x"7e", -- $08293
          33428 => x"7e", -- $08294
          33429 => x"7f", -- $08295
          33430 => x"7f", -- $08296
          33431 => x"7f", -- $08297
          33432 => x"7f", -- $08298
          33433 => x"7f", -- $08299
          33434 => x"7f", -- $0829a
          33435 => x"7f", -- $0829b
          33436 => x"7f", -- $0829c
          33437 => x"7f", -- $0829d
          33438 => x"7e", -- $0829e
          33439 => x"7e", -- $0829f
          33440 => x"7e", -- $082a0
          33441 => x"7e", -- $082a1
          33442 => x"7e", -- $082a2
          33443 => x"7e", -- $082a3
          33444 => x"7e", -- $082a4
          33445 => x"7e", -- $082a5
          33446 => x"7e", -- $082a6
          33447 => x"7e", -- $082a7
          33448 => x"7e", -- $082a8
          33449 => x"7e", -- $082a9
          33450 => x"7e", -- $082aa
          33451 => x"7e", -- $082ab
          33452 => x"7d", -- $082ac
          33453 => x"7d", -- $082ad
          33454 => x"7e", -- $082ae
          33455 => x"7e", -- $082af
          33456 => x"7e", -- $082b0
          33457 => x"7e", -- $082b1
          33458 => x"7e", -- $082b2
          33459 => x"7e", -- $082b3
          33460 => x"7e", -- $082b4
          33461 => x"7e", -- $082b5
          33462 => x"7e", -- $082b6
          33463 => x"7e", -- $082b7
          33464 => x"7e", -- $082b8
          33465 => x"7e", -- $082b9
          33466 => x"7e", -- $082ba
          33467 => x"7e", -- $082bb
          33468 => x"7e", -- $082bc
          33469 => x"7e", -- $082bd
          33470 => x"7e", -- $082be
          33471 => x"7e", -- $082bf
          33472 => x"7e", -- $082c0
          33473 => x"7e", -- $082c1
          33474 => x"7e", -- $082c2
          33475 => x"7e", -- $082c3
          33476 => x"7e", -- $082c4
          33477 => x"7e", -- $082c5
          33478 => x"7e", -- $082c6
          33479 => x"7e", -- $082c7
          33480 => x"7e", -- $082c8
          33481 => x"7d", -- $082c9
          33482 => x"7d", -- $082ca
          33483 => x"7d", -- $082cb
          33484 => x"7d", -- $082cc
          33485 => x"7d", -- $082cd
          33486 => x"7d", -- $082ce
          33487 => x"7d", -- $082cf
          33488 => x"7d", -- $082d0
          33489 => x"7d", -- $082d1
          33490 => x"7d", -- $082d2
          33491 => x"7e", -- $082d3
          33492 => x"7e", -- $082d4
          33493 => x"7e", -- $082d5
          33494 => x"7e", -- $082d6
          33495 => x"7e", -- $082d7
          33496 => x"7e", -- $082d8
          33497 => x"7e", -- $082d9
          33498 => x"7f", -- $082da
          33499 => x"7f", -- $082db
          33500 => x"7f", -- $082dc
          33501 => x"7f", -- $082dd
          33502 => x"7f", -- $082de
          33503 => x"7f", -- $082df
          33504 => x"7f", -- $082e0
          33505 => x"7f", -- $082e1
          33506 => x"7f", -- $082e2
          33507 => x"7e", -- $082e3
          33508 => x"7e", -- $082e4
          33509 => x"7e", -- $082e5
          33510 => x"7e", -- $082e6
          33511 => x"7e", -- $082e7
          33512 => x"7e", -- $082e8
          33513 => x"7e", -- $082e9
          33514 => x"7e", -- $082ea
          33515 => x"7e", -- $082eb
          33516 => x"7e", -- $082ec
          33517 => x"7e", -- $082ed
          33518 => x"7e", -- $082ee
          33519 => x"7e", -- $082ef
          33520 => x"7e", -- $082f0
          33521 => x"7e", -- $082f1
          33522 => x"7e", -- $082f2
          33523 => x"7e", -- $082f3
          33524 => x"7f", -- $082f4
          33525 => x"7f", -- $082f5
          33526 => x"7f", -- $082f6
          33527 => x"7f", -- $082f7
          33528 => x"7f", -- $082f8
          33529 => x"7f", -- $082f9
          33530 => x"7f", -- $082fa
          33531 => x"7f", -- $082fb
          33532 => x"7f", -- $082fc
          33533 => x"7f", -- $082fd
          33534 => x"7f", -- $082fe
          33535 => x"7f", -- $082ff
          33536 => x"7f", -- $08300
          33537 => x"7f", -- $08301
          33538 => x"7f", -- $08302
          33539 => x"7f", -- $08303
          33540 => x"7f", -- $08304
          33541 => x"7f", -- $08305
          33542 => x"7f", -- $08306
          33543 => x"7f", -- $08307
          33544 => x"7f", -- $08308
          33545 => x"7e", -- $08309
          33546 => x"7e", -- $0830a
          33547 => x"7e", -- $0830b
          33548 => x"7e", -- $0830c
          33549 => x"7e", -- $0830d
          33550 => x"7e", -- $0830e
          33551 => x"7e", -- $0830f
          33552 => x"7e", -- $08310
          33553 => x"7e", -- $08311
          33554 => x"7e", -- $08312
          33555 => x"7e", -- $08313
          33556 => x"7f", -- $08314
          33557 => x"7f", -- $08315
          33558 => x"7f", -- $08316
          33559 => x"7f", -- $08317
          33560 => x"7f", -- $08318
          33561 => x"7f", -- $08319
          33562 => x"7f", -- $0831a
          33563 => x"7f", -- $0831b
          33564 => x"7f", -- $0831c
          33565 => x"7f", -- $0831d
          33566 => x"7f", -- $0831e
          33567 => x"7f", -- $0831f
          33568 => x"7f", -- $08320
          33569 => x"7f", -- $08321
          33570 => x"7f", -- $08322
          33571 => x"7f", -- $08323
          33572 => x"7f", -- $08324
          33573 => x"7f", -- $08325
          33574 => x"7f", -- $08326
          33575 => x"7f", -- $08327
          33576 => x"7f", -- $08328
          33577 => x"7e", -- $08329
          33578 => x"7e", -- $0832a
          33579 => x"7e", -- $0832b
          33580 => x"7e", -- $0832c
          33581 => x"7e", -- $0832d
          33582 => x"7e", -- $0832e
          33583 => x"7e", -- $0832f
          33584 => x"7e", -- $08330
          33585 => x"7e", -- $08331
          33586 => x"7e", -- $08332
          33587 => x"7e", -- $08333
          33588 => x"7f", -- $08334
          33589 => x"7f", -- $08335
          33590 => x"7f", -- $08336
          33591 => x"7f", -- $08337
          33592 => x"7f", -- $08338
          33593 => x"7f", -- $08339
          33594 => x"7f", -- $0833a
          33595 => x"7f", -- $0833b
          33596 => x"7f", -- $0833c
          33597 => x"7f", -- $0833d
          33598 => x"7f", -- $0833e
          33599 => x"7f", -- $0833f
          33600 => x"7f", -- $08340
          33601 => x"7f", -- $08341
          33602 => x"7f", -- $08342
          33603 => x"7f", -- $08343
          33604 => x"7f", -- $08344
          33605 => x"7f", -- $08345
          33606 => x"7f", -- $08346
          33607 => x"7e", -- $08347
          33608 => x"7e", -- $08348
          33609 => x"7e", -- $08349
          33610 => x"7e", -- $0834a
          33611 => x"7e", -- $0834b
          33612 => x"7e", -- $0834c
          33613 => x"7e", -- $0834d
          33614 => x"7e", -- $0834e
          33615 => x"7e", -- $0834f
          33616 => x"7e", -- $08350
          33617 => x"7e", -- $08351
          33618 => x"7e", -- $08352
          33619 => x"7f", -- $08353
          33620 => x"7f", -- $08354
          33621 => x"7f", -- $08355
          33622 => x"7f", -- $08356
          33623 => x"7f", -- $08357
          33624 => x"7f", -- $08358
          33625 => x"7f", -- $08359
          33626 => x"80", -- $0835a
          33627 => x"80", -- $0835b
          33628 => x"80", -- $0835c
          33629 => x"80", -- $0835d
          33630 => x"80", -- $0835e
          33631 => x"80", -- $0835f
          33632 => x"7f", -- $08360
          33633 => x"7f", -- $08361
          33634 => x"7f", -- $08362
          33635 => x"7f", -- $08363
          33636 => x"7f", -- $08364
          33637 => x"7f", -- $08365
          33638 => x"7f", -- $08366
          33639 => x"7f", -- $08367
          33640 => x"7f", -- $08368
          33641 => x"7f", -- $08369
          33642 => x"7f", -- $0836a
          33643 => x"7f", -- $0836b
          33644 => x"7e", -- $0836c
          33645 => x"7e", -- $0836d
          33646 => x"7e", -- $0836e
          33647 => x"7e", -- $0836f
          33648 => x"7f", -- $08370
          33649 => x"7f", -- $08371
          33650 => x"7f", -- $08372
          33651 => x"7f", -- $08373
          33652 => x"7f", -- $08374
          33653 => x"80", -- $08375
          33654 => x"80", -- $08376
          33655 => x"80", -- $08377
          33656 => x"80", -- $08378
          33657 => x"80", -- $08379
          33658 => x"80", -- $0837a
          33659 => x"80", -- $0837b
          33660 => x"80", -- $0837c
          33661 => x"80", -- $0837d
          33662 => x"80", -- $0837e
          33663 => x"80", -- $0837f
          33664 => x"80", -- $08380
          33665 => x"80", -- $08381
          33666 => x"80", -- $08382
          33667 => x"80", -- $08383
          33668 => x"80", -- $08384
          33669 => x"80", -- $08385
          33670 => x"80", -- $08386
          33671 => x"80", -- $08387
          33672 => x"7f", -- $08388
          33673 => x"7f", -- $08389
          33674 => x"7f", -- $0838a
          33675 => x"7f", -- $0838b
          33676 => x"7f", -- $0838c
          33677 => x"7f", -- $0838d
          33678 => x"7f", -- $0838e
          33679 => x"80", -- $0838f
          33680 => x"80", -- $08390
          33681 => x"80", -- $08391
          33682 => x"80", -- $08392
          33683 => x"80", -- $08393
          33684 => x"80", -- $08394
          33685 => x"80", -- $08395
          33686 => x"80", -- $08396
          33687 => x"80", -- $08397
          33688 => x"80", -- $08398
          33689 => x"80", -- $08399
          33690 => x"81", -- $0839a
          33691 => x"81", -- $0839b
          33692 => x"81", -- $0839c
          33693 => x"81", -- $0839d
          33694 => x"81", -- $0839e
          33695 => x"81", -- $0839f
          33696 => x"81", -- $083a0
          33697 => x"81", -- $083a1
          33698 => x"80", -- $083a2
          33699 => x"80", -- $083a3
          33700 => x"80", -- $083a4
          33701 => x"80", -- $083a5
          33702 => x"80", -- $083a6
          33703 => x"80", -- $083a7
          33704 => x"80", -- $083a8
          33705 => x"80", -- $083a9
          33706 => x"80", -- $083aa
          33707 => x"80", -- $083ab
          33708 => x"80", -- $083ac
          33709 => x"80", -- $083ad
          33710 => x"80", -- $083ae
          33711 => x"80", -- $083af
          33712 => x"80", -- $083b0
          33713 => x"80", -- $083b1
          33714 => x"80", -- $083b2
          33715 => x"80", -- $083b3
          33716 => x"81", -- $083b4
          33717 => x"81", -- $083b5
          33718 => x"81", -- $083b6
          33719 => x"81", -- $083b7
          33720 => x"82", -- $083b8
          33721 => x"81", -- $083b9
          33722 => x"82", -- $083ba
          33723 => x"82", -- $083bb
          33724 => x"82", -- $083bc
          33725 => x"82", -- $083bd
          33726 => x"81", -- $083be
          33727 => x"81", -- $083bf
          33728 => x"81", -- $083c0
          33729 => x"81", -- $083c1
          33730 => x"81", -- $083c2
          33731 => x"81", -- $083c3
          33732 => x"81", -- $083c4
          33733 => x"81", -- $083c5
          33734 => x"81", -- $083c6
          33735 => x"80", -- $083c7
          33736 => x"80", -- $083c8
          33737 => x"80", -- $083c9
          33738 => x"80", -- $083ca
          33739 => x"80", -- $083cb
          33740 => x"80", -- $083cc
          33741 => x"80", -- $083cd
          33742 => x"80", -- $083ce
          33743 => x"80", -- $083cf
          33744 => x"81", -- $083d0
          33745 => x"81", -- $083d1
          33746 => x"81", -- $083d2
          33747 => x"81", -- $083d3
          33748 => x"81", -- $083d4
          33749 => x"81", -- $083d5
          33750 => x"82", -- $083d6
          33751 => x"82", -- $083d7
          33752 => x"82", -- $083d8
          33753 => x"82", -- $083d9
          33754 => x"82", -- $083da
          33755 => x"82", -- $083db
          33756 => x"82", -- $083dc
          33757 => x"82", -- $083dd
          33758 => x"82", -- $083de
          33759 => x"82", -- $083df
          33760 => x"82", -- $083e0
          33761 => x"81", -- $083e1
          33762 => x"81", -- $083e2
          33763 => x"81", -- $083e3
          33764 => x"81", -- $083e4
          33765 => x"81", -- $083e5
          33766 => x"81", -- $083e6
          33767 => x"81", -- $083e7
          33768 => x"81", -- $083e8
          33769 => x"81", -- $083e9
          33770 => x"80", -- $083ea
          33771 => x"81", -- $083eb
          33772 => x"81", -- $083ec
          33773 => x"80", -- $083ed
          33774 => x"80", -- $083ee
          33775 => x"81", -- $083ef
          33776 => x"81", -- $083f0
          33777 => x"81", -- $083f1
          33778 => x"81", -- $083f2
          33779 => x"81", -- $083f3
          33780 => x"81", -- $083f4
          33781 => x"81", -- $083f5
          33782 => x"82", -- $083f6
          33783 => x"82", -- $083f7
          33784 => x"82", -- $083f8
          33785 => x"82", -- $083f9
          33786 => x"82", -- $083fa
          33787 => x"82", -- $083fb
          33788 => x"82", -- $083fc
          33789 => x"82", -- $083fd
          33790 => x"81", -- $083fe
          33791 => x"81", -- $083ff
          33792 => x"81", -- $08400
          33793 => x"81", -- $08401
          33794 => x"81", -- $08402
          33795 => x"81", -- $08403
          33796 => x"81", -- $08404
          33797 => x"81", -- $08405
          33798 => x"80", -- $08406
          33799 => x"80", -- $08407
          33800 => x"80", -- $08408
          33801 => x"80", -- $08409
          33802 => x"80", -- $0840a
          33803 => x"80", -- $0840b
          33804 => x"80", -- $0840c
          33805 => x"80", -- $0840d
          33806 => x"81", -- $0840e
          33807 => x"81", -- $0840f
          33808 => x"81", -- $08410
          33809 => x"81", -- $08411
          33810 => x"81", -- $08412
          33811 => x"81", -- $08413
          33812 => x"81", -- $08414
          33813 => x"81", -- $08415
          33814 => x"81", -- $08416
          33815 => x"81", -- $08417
          33816 => x"82", -- $08418
          33817 => x"82", -- $08419
          33818 => x"82", -- $0841a
          33819 => x"82", -- $0841b
          33820 => x"82", -- $0841c
          33821 => x"82", -- $0841d
          33822 => x"82", -- $0841e
          33823 => x"82", -- $0841f
          33824 => x"81", -- $08420
          33825 => x"81", -- $08421
          33826 => x"81", -- $08422
          33827 => x"81", -- $08423
          33828 => x"81", -- $08424
          33829 => x"81", -- $08425
          33830 => x"81", -- $08426
          33831 => x"81", -- $08427
          33832 => x"81", -- $08428
          33833 => x"81", -- $08429
          33834 => x"81", -- $0842a
          33835 => x"81", -- $0842b
          33836 => x"81", -- $0842c
          33837 => x"81", -- $0842d
          33838 => x"81", -- $0842e
          33839 => x"81", -- $0842f
          33840 => x"81", -- $08430
          33841 => x"82", -- $08431
          33842 => x"82", -- $08432
          33843 => x"82", -- $08433
          33844 => x"82", -- $08434
          33845 => x"82", -- $08435
          33846 => x"82", -- $08436
          33847 => x"82", -- $08437
          33848 => x"82", -- $08438
          33849 => x"82", -- $08439
          33850 => x"82", -- $0843a
          33851 => x"82", -- $0843b
          33852 => x"82", -- $0843c
          33853 => x"82", -- $0843d
          33854 => x"82", -- $0843e
          33855 => x"82", -- $0843f
          33856 => x"82", -- $08440
          33857 => x"82", -- $08441
          33858 => x"82", -- $08442
          33859 => x"81", -- $08443
          33860 => x"81", -- $08444
          33861 => x"81", -- $08445
          33862 => x"81", -- $08446
          33863 => x"81", -- $08447
          33864 => x"81", -- $08448
          33865 => x"81", -- $08449
          33866 => x"81", -- $0844a
          33867 => x"81", -- $0844b
          33868 => x"81", -- $0844c
          33869 => x"81", -- $0844d
          33870 => x"82", -- $0844e
          33871 => x"82", -- $0844f
          33872 => x"82", -- $08450
          33873 => x"82", -- $08451
          33874 => x"82", -- $08452
          33875 => x"82", -- $08453
          33876 => x"82", -- $08454
          33877 => x"82", -- $08455
          33878 => x"82", -- $08456
          33879 => x"82", -- $08457
          33880 => x"82", -- $08458
          33881 => x"82", -- $08459
          33882 => x"82", -- $0845a
          33883 => x"82", -- $0845b
          33884 => x"82", -- $0845c
          33885 => x"82", -- $0845d
          33886 => x"82", -- $0845e
          33887 => x"82", -- $0845f
          33888 => x"82", -- $08460
          33889 => x"82", -- $08461
          33890 => x"82", -- $08462
          33891 => x"82", -- $08463
          33892 => x"82", -- $08464
          33893 => x"81", -- $08465
          33894 => x"81", -- $08466
          33895 => x"81", -- $08467
          33896 => x"81", -- $08468
          33897 => x"81", -- $08469
          33898 => x"81", -- $0846a
          33899 => x"81", -- $0846b
          33900 => x"81", -- $0846c
          33901 => x"82", -- $0846d
          33902 => x"82", -- $0846e
          33903 => x"82", -- $0846f
          33904 => x"82", -- $08470
          33905 => x"82", -- $08471
          33906 => x"82", -- $08472
          33907 => x"82", -- $08473
          33908 => x"82", -- $08474
          33909 => x"82", -- $08475
          33910 => x"82", -- $08476
          33911 => x"82", -- $08477
          33912 => x"82", -- $08478
          33913 => x"82", -- $08479
          33914 => x"82", -- $0847a
          33915 => x"82", -- $0847b
          33916 => x"82", -- $0847c
          33917 => x"82", -- $0847d
          33918 => x"82", -- $0847e
          33919 => x"82", -- $0847f
          33920 => x"82", -- $08480
          33921 => x"81", -- $08481
          33922 => x"81", -- $08482
          33923 => x"81", -- $08483
          33924 => x"81", -- $08484
          33925 => x"81", -- $08485
          33926 => x"81", -- $08486
          33927 => x"81", -- $08487
          33928 => x"81", -- $08488
          33929 => x"81", -- $08489
          33930 => x"81", -- $0848a
          33931 => x"81", -- $0848b
          33932 => x"82", -- $0848c
          33933 => x"82", -- $0848d
          33934 => x"82", -- $0848e
          33935 => x"82", -- $0848f
          33936 => x"82", -- $08490
          33937 => x"82", -- $08491
          33938 => x"82", -- $08492
          33939 => x"82", -- $08493
          33940 => x"82", -- $08494
          33941 => x"82", -- $08495
          33942 => x"82", -- $08496
          33943 => x"82", -- $08497
          33944 => x"82", -- $08498
          33945 => x"82", -- $08499
          33946 => x"82", -- $0849a
          33947 => x"82", -- $0849b
          33948 => x"82", -- $0849c
          33949 => x"82", -- $0849d
          33950 => x"82", -- $0849e
          33951 => x"82", -- $0849f
          33952 => x"82", -- $084a0
          33953 => x"82", -- $084a1
          33954 => x"81", -- $084a2
          33955 => x"81", -- $084a3
          33956 => x"81", -- $084a4
          33957 => x"81", -- $084a5
          33958 => x"81", -- $084a6
          33959 => x"81", -- $084a7
          33960 => x"81", -- $084a8
          33961 => x"81", -- $084a9
          33962 => x"81", -- $084aa
          33963 => x"81", -- $084ab
          33964 => x"81", -- $084ac
          33965 => x"81", -- $084ad
          33966 => x"81", -- $084ae
          33967 => x"81", -- $084af
          33968 => x"81", -- $084b0
          33969 => x"81", -- $084b1
          33970 => x"81", -- $084b2
          33971 => x"81", -- $084b3
          33972 => x"81", -- $084b4
          33973 => x"81", -- $084b5
          33974 => x"81", -- $084b6
          33975 => x"81", -- $084b7
          33976 => x"81", -- $084b8
          33977 => x"81", -- $084b9
          33978 => x"81", -- $084ba
          33979 => x"81", -- $084bb
          33980 => x"81", -- $084bc
          33981 => x"81", -- $084bd
          33982 => x"81", -- $084be
          33983 => x"81", -- $084bf
          33984 => x"81", -- $084c0
          33985 => x"81", -- $084c1
          33986 => x"81", -- $084c2
          33987 => x"81", -- $084c3
          33988 => x"81", -- $084c4
          33989 => x"81", -- $084c5
          33990 => x"81", -- $084c6
          33991 => x"81", -- $084c7
          33992 => x"81", -- $084c8
          33993 => x"81", -- $084c9
          33994 => x"81", -- $084ca
          33995 => x"81", -- $084cb
          33996 => x"81", -- $084cc
          33997 => x"81", -- $084cd
          33998 => x"81", -- $084ce
          33999 => x"81", -- $084cf
          34000 => x"81", -- $084d0
          34001 => x"81", -- $084d1
          34002 => x"81", -- $084d2
          34003 => x"81", -- $084d3
          34004 => x"81", -- $084d4
          34005 => x"81", -- $084d5
          34006 => x"81", -- $084d6
          34007 => x"81", -- $084d7
          34008 => x"81", -- $084d8
          34009 => x"81", -- $084d9
          34010 => x"81", -- $084da
          34011 => x"81", -- $084db
          34012 => x"81", -- $084dc
          34013 => x"81", -- $084dd
          34014 => x"81", -- $084de
          34015 => x"81", -- $084df
          34016 => x"81", -- $084e0
          34017 => x"80", -- $084e1
          34018 => x"80", -- $084e2
          34019 => x"80", -- $084e3
          34020 => x"80", -- $084e4
          34021 => x"80", -- $084e5
          34022 => x"80", -- $084e6
          34023 => x"80", -- $084e7
          34024 => x"80", -- $084e8
          34025 => x"80", -- $084e9
          34026 => x"80", -- $084ea
          34027 => x"80", -- $084eb
          34028 => x"80", -- $084ec
          34029 => x"80", -- $084ed
          34030 => x"80", -- $084ee
          34031 => x"80", -- $084ef
          34032 => x"80", -- $084f0
          34033 => x"80", -- $084f1
          34034 => x"80", -- $084f2
          34035 => x"80", -- $084f3
          34036 => x"80", -- $084f4
          34037 => x"80", -- $084f5
          34038 => x"80", -- $084f6
          34039 => x"80", -- $084f7
          34040 => x"80", -- $084f8
          34041 => x"80", -- $084f9
          34042 => x"80", -- $084fa
          34043 => x"80", -- $084fb
          34044 => x"80", -- $084fc
          34045 => x"80", -- $084fd
          34046 => x"80", -- $084fe
          34047 => x"80", -- $084ff
          34048 => x"80", -- $08500
          34049 => x"80", -- $08501
          34050 => x"80", -- $08502
          34051 => x"80", -- $08503
          34052 => x"80", -- $08504
          34053 => x"80", -- $08505
          34054 => x"80", -- $08506
          34055 => x"80", -- $08507
          34056 => x"80", -- $08508
          34057 => x"80", -- $08509
          34058 => x"80", -- $0850a
          34059 => x"80", -- $0850b
          34060 => x"80", -- $0850c
          34061 => x"80", -- $0850d
          34062 => x"80", -- $0850e
          34063 => x"80", -- $0850f
          34064 => x"80", -- $08510
          34065 => x"80", -- $08511
          34066 => x"80", -- $08512
          34067 => x"80", -- $08513
          34068 => x"80", -- $08514
          34069 => x"80", -- $08515
          34070 => x"80", -- $08516
          34071 => x"80", -- $08517
          34072 => x"80", -- $08518
          34073 => x"80", -- $08519
          34074 => x"80", -- $0851a
          34075 => x"80", -- $0851b
          34076 => x"80", -- $0851c
          34077 => x"80", -- $0851d
          34078 => x"80", -- $0851e
          34079 => x"80", -- $0851f
          34080 => x"80", -- $08520
          34081 => x"80", -- $08521
          34082 => x"80", -- $08522
          34083 => x"80", -- $08523
          34084 => x"80", -- $08524
          34085 => x"80", -- $08525
          34086 => x"80", -- $08526
          34087 => x"80", -- $08527
          34088 => x"80", -- $08528
          34089 => x"7f", -- $08529
          34090 => x"7f", -- $0852a
          34091 => x"7f", -- $0852b
          34092 => x"7f", -- $0852c
          34093 => x"7f", -- $0852d
          34094 => x"80", -- $0852e
          34095 => x"80", -- $0852f
          34096 => x"80", -- $08530
          34097 => x"80", -- $08531
          34098 => x"80", -- $08532
          34099 => x"80", -- $08533
          34100 => x"80", -- $08534
          34101 => x"80", -- $08535
          34102 => x"80", -- $08536
          34103 => x"80", -- $08537
          34104 => x"80", -- $08538
          34105 => x"80", -- $08539
          34106 => x"80", -- $0853a
          34107 => x"80", -- $0853b
          34108 => x"80", -- $0853c
          34109 => x"80", -- $0853d
          34110 => x"80", -- $0853e
          34111 => x"80", -- $0853f
          34112 => x"80", -- $08540
          34113 => x"7f", -- $08541
          34114 => x"7f", -- $08542
          34115 => x"7f", -- $08543
          34116 => x"7f", -- $08544
          34117 => x"7f", -- $08545
          34118 => x"7f", -- $08546
          34119 => x"7f", -- $08547
          34120 => x"7f", -- $08548
          34121 => x"7f", -- $08549
          34122 => x"7f", -- $0854a
          34123 => x"7f", -- $0854b
          34124 => x"7f", -- $0854c
          34125 => x"7f", -- $0854d
          34126 => x"7f", -- $0854e
          34127 => x"80", -- $0854f
          34128 => x"7f", -- $08550
          34129 => x"80", -- $08551
          34130 => x"80", -- $08552
          34131 => x"80", -- $08553
          34132 => x"80", -- $08554
          34133 => x"80", -- $08555
          34134 => x"80", -- $08556
          34135 => x"80", -- $08557
          34136 => x"80", -- $08558
          34137 => x"80", -- $08559
          34138 => x"80", -- $0855a
          34139 => x"80", -- $0855b
          34140 => x"80", -- $0855c
          34141 => x"80", -- $0855d
          34142 => x"80", -- $0855e
          34143 => x"7f", -- $0855f
          34144 => x"7f", -- $08560
          34145 => x"7f", -- $08561
          34146 => x"7f", -- $08562
          34147 => x"7f", -- $08563
          34148 => x"80", -- $08564
          34149 => x"7f", -- $08565
          34150 => x"7f", -- $08566
          34151 => x"80", -- $08567
          34152 => x"7f", -- $08568
          34153 => x"80", -- $08569
          34154 => x"7f", -- $0856a
          34155 => x"7f", -- $0856b
          34156 => x"7f", -- $0856c
          34157 => x"7f", -- $0856d
          34158 => x"7f", -- $0856e
          34159 => x"7f", -- $0856f
          34160 => x"7f", -- $08570
          34161 => x"7f", -- $08571
          34162 => x"7f", -- $08572
          34163 => x"80", -- $08573
          34164 => x"80", -- $08574
          34165 => x"7f", -- $08575
          34166 => x"7f", -- $08576
          34167 => x"7f", -- $08577
          34168 => x"7f", -- $08578
          34169 => x"7f", -- $08579
          34170 => x"7f", -- $0857a
          34171 => x"7f", -- $0857b
          34172 => x"7f", -- $0857c
          34173 => x"7f", -- $0857d
          34174 => x"7f", -- $0857e
          34175 => x"7f", -- $0857f
          34176 => x"7f", -- $08580
          34177 => x"7f", -- $08581
          34178 => x"7f", -- $08582
          34179 => x"7f", -- $08583
          34180 => x"7f", -- $08584
          34181 => x"7f", -- $08585
          34182 => x"7f", -- $08586
          34183 => x"7f", -- $08587
          34184 => x"7f", -- $08588
          34185 => x"7f", -- $08589
          34186 => x"7f", -- $0858a
          34187 => x"7f", -- $0858b
          34188 => x"7f", -- $0858c
          34189 => x"7f", -- $0858d
          34190 => x"7f", -- $0858e
          34191 => x"7f", -- $0858f
          34192 => x"7f", -- $08590
          34193 => x"7f", -- $08591
          34194 => x"7f", -- $08592
          34195 => x"7f", -- $08593
          34196 => x"7f", -- $08594
          34197 => x"7f", -- $08595
          34198 => x"7f", -- $08596
          34199 => x"7f", -- $08597
          34200 => x"7f", -- $08598
          34201 => x"7f", -- $08599
          34202 => x"7f", -- $0859a
          34203 => x"7f", -- $0859b
          34204 => x"7e", -- $0859c
          34205 => x"7e", -- $0859d
          34206 => x"7e", -- $0859e
          34207 => x"7e", -- $0859f
          34208 => x"7e", -- $085a0
          34209 => x"7e", -- $085a1
          34210 => x"7e", -- $085a2
          34211 => x"7e", -- $085a3
          34212 => x"7e", -- $085a4
          34213 => x"7e", -- $085a5
          34214 => x"7e", -- $085a6
          34215 => x"7e", -- $085a7
          34216 => x"7e", -- $085a8
          34217 => x"7e", -- $085a9
          34218 => x"7e", -- $085aa
          34219 => x"7e", -- $085ab
          34220 => x"7e", -- $085ac
          34221 => x"7e", -- $085ad
          34222 => x"7e", -- $085ae
          34223 => x"7e", -- $085af
          34224 => x"7e", -- $085b0
          34225 => x"7e", -- $085b1
          34226 => x"7e", -- $085b2
          34227 => x"7e", -- $085b3
          34228 => x"7e", -- $085b4
          34229 => x"7e", -- $085b5
          34230 => x"7e", -- $085b6
          34231 => x"7e", -- $085b7
          34232 => x"7e", -- $085b8
          34233 => x"7e", -- $085b9
          34234 => x"7e", -- $085ba
          34235 => x"7e", -- $085bb
          34236 => x"7e", -- $085bc
          34237 => x"7e", -- $085bd
          34238 => x"7e", -- $085be
          34239 => x"7e", -- $085bf
          34240 => x"7e", -- $085c0
          34241 => x"7e", -- $085c1
          34242 => x"7e", -- $085c2
          34243 => x"7e", -- $085c3
          34244 => x"7e", -- $085c4
          34245 => x"7e", -- $085c5
          34246 => x"7e", -- $085c6
          34247 => x"7e", -- $085c7
          34248 => x"7e", -- $085c8
          34249 => x"7e", -- $085c9
          34250 => x"7e", -- $085ca
          34251 => x"7e", -- $085cb
          34252 => x"7e", -- $085cc
          34253 => x"7e", -- $085cd
          34254 => x"7e", -- $085ce
          34255 => x"7e", -- $085cf
          34256 => x"7e", -- $085d0
          34257 => x"7e", -- $085d1
          34258 => x"7d", -- $085d2
          34259 => x"7d", -- $085d3
          34260 => x"7d", -- $085d4
          34261 => x"7d", -- $085d5
          34262 => x"7d", -- $085d6
          34263 => x"7d", -- $085d7
          34264 => x"7d", -- $085d8
          34265 => x"7d", -- $085d9
          34266 => x"7e", -- $085da
          34267 => x"7e", -- $085db
          34268 => x"7e", -- $085dc
          34269 => x"7e", -- $085dd
          34270 => x"7e", -- $085de
          34271 => x"7e", -- $085df
          34272 => x"7e", -- $085e0
          34273 => x"7e", -- $085e1
          34274 => x"7e", -- $085e2
          34275 => x"7e", -- $085e3
          34276 => x"7e", -- $085e4
          34277 => x"7e", -- $085e5
          34278 => x"7e", -- $085e6
          34279 => x"7e", -- $085e7
          34280 => x"7e", -- $085e8
          34281 => x"7e", -- $085e9
          34282 => x"7e", -- $085ea
          34283 => x"7e", -- $085eb
          34284 => x"7e", -- $085ec
          34285 => x"7e", -- $085ed
          34286 => x"7e", -- $085ee
          34287 => x"7e", -- $085ef
          34288 => x"7e", -- $085f0
          34289 => x"7e", -- $085f1
          34290 => x"7e", -- $085f2
          34291 => x"7e", -- $085f3
          34292 => x"7e", -- $085f4
          34293 => x"7e", -- $085f5
          34294 => x"7e", -- $085f6
          34295 => x"7e", -- $085f7
          34296 => x"7e", -- $085f8
          34297 => x"7e", -- $085f9
          34298 => x"7e", -- $085fa
          34299 => x"7e", -- $085fb
          34300 => x"7e", -- $085fc
          34301 => x"7f", -- $085fd
          34302 => x"7f", -- $085fe
          34303 => x"7f", -- $085ff
          34304 => x"7f", -- $08600
          34305 => x"7f", -- $08601
          34306 => x"7f", -- $08602
          34307 => x"7f", -- $08603
          34308 => x"7f", -- $08604
          34309 => x"7f", -- $08605
          34310 => x"7f", -- $08606
          34311 => x"7f", -- $08607
          34312 => x"7f", -- $08608
          34313 => x"7f", -- $08609
          34314 => x"7f", -- $0860a
          34315 => x"7f", -- $0860b
          34316 => x"7f", -- $0860c
          34317 => x"7f", -- $0860d
          34318 => x"7f", -- $0860e
          34319 => x"7f", -- $0860f
          34320 => x"7f", -- $08610
          34321 => x"7f", -- $08611
          34322 => x"7f", -- $08612
          34323 => x"7f", -- $08613
          34324 => x"7f", -- $08614
          34325 => x"7f", -- $08615
          34326 => x"7f", -- $08616
          34327 => x"7f", -- $08617
          34328 => x"7f", -- $08618
          34329 => x"7f", -- $08619
          34330 => x"7f", -- $0861a
          34331 => x"7f", -- $0861b
          34332 => x"7f", -- $0861c
          34333 => x"7f", -- $0861d
          34334 => x"80", -- $0861e
          34335 => x"80", -- $0861f
          34336 => x"7f", -- $08620
          34337 => x"80", -- $08621
          34338 => x"80", -- $08622
          34339 => x"80", -- $08623
          34340 => x"80", -- $08624
          34341 => x"80", -- $08625
          34342 => x"80", -- $08626
          34343 => x"80", -- $08627
          34344 => x"80", -- $08628
          34345 => x"80", -- $08629
          34346 => x"80", -- $0862a
          34347 => x"80", -- $0862b
          34348 => x"80", -- $0862c
          34349 => x"7f", -- $0862d
          34350 => x"7f", -- $0862e
          34351 => x"7f", -- $0862f
          34352 => x"7f", -- $08630
          34353 => x"7f", -- $08631
          34354 => x"7f", -- $08632
          34355 => x"7f", -- $08633
          34356 => x"7f", -- $08634
          34357 => x"7f", -- $08635
          34358 => x"7f", -- $08636
          34359 => x"7f", -- $08637
          34360 => x"7f", -- $08638
          34361 => x"80", -- $08639
          34362 => x"80", -- $0863a
          34363 => x"80", -- $0863b
          34364 => x"80", -- $0863c
          34365 => x"80", -- $0863d
          34366 => x"80", -- $0863e
          34367 => x"80", -- $0863f
          34368 => x"80", -- $08640
          34369 => x"80", -- $08641
          34370 => x"80", -- $08642
          34371 => x"80", -- $08643
          34372 => x"80", -- $08644
          34373 => x"80", -- $08645
          34374 => x"80", -- $08646
          34375 => x"80", -- $08647
          34376 => x"80", -- $08648
          34377 => x"80", -- $08649
          34378 => x"80", -- $0864a
          34379 => x"80", -- $0864b
          34380 => x"80", -- $0864c
          34381 => x"80", -- $0864d
          34382 => x"80", -- $0864e
          34383 => x"80", -- $0864f
          34384 => x"80", -- $08650
          34385 => x"80", -- $08651
          34386 => x"80", -- $08652
          34387 => x"7f", -- $08653
          34388 => x"7f", -- $08654
          34389 => x"7f", -- $08655
          34390 => x"7f", -- $08656
          34391 => x"80", -- $08657
          34392 => x"80", -- $08658
          34393 => x"80", -- $08659
          34394 => x"80", -- $0865a
          34395 => x"80", -- $0865b
          34396 => x"80", -- $0865c
          34397 => x"80", -- $0865d
          34398 => x"80", -- $0865e
          34399 => x"80", -- $0865f
          34400 => x"80", -- $08660
          34401 => x"80", -- $08661
          34402 => x"80", -- $08662
          34403 => x"80", -- $08663
          34404 => x"80", -- $08664
          34405 => x"80", -- $08665
          34406 => x"80", -- $08666
          34407 => x"80", -- $08667
          34408 => x"80", -- $08668
          34409 => x"80", -- $08669
          34410 => x"80", -- $0866a
          34411 => x"80", -- $0866b
          34412 => x"80", -- $0866c
          34413 => x"80", -- $0866d
          34414 => x"80", -- $0866e
          34415 => x"80", -- $0866f
          34416 => x"80", -- $08670
          34417 => x"80", -- $08671
          34418 => x"80", -- $08672
          34419 => x"80", -- $08673
          34420 => x"80", -- $08674
          34421 => x"80", -- $08675
          34422 => x"80", -- $08676
          34423 => x"80", -- $08677
          34424 => x"80", -- $08678
          34425 => x"80", -- $08679
          34426 => x"80", -- $0867a
          34427 => x"80", -- $0867b
          34428 => x"80", -- $0867c
          34429 => x"80", -- $0867d
          34430 => x"80", -- $0867e
          34431 => x"80", -- $0867f
          34432 => x"80", -- $08680
          34433 => x"80", -- $08681
          34434 => x"80", -- $08682
          34435 => x"80", -- $08683
          34436 => x"80", -- $08684
          34437 => x"80", -- $08685
          34438 => x"80", -- $08686
          34439 => x"80", -- $08687
          34440 => x"80", -- $08688
          34441 => x"80", -- $08689
          34442 => x"80", -- $0868a
          34443 => x"80", -- $0868b
          34444 => x"80", -- $0868c
          34445 => x"80", -- $0868d
          34446 => x"80", -- $0868e
          34447 => x"80", -- $0868f
          34448 => x"80", -- $08690
          34449 => x"80", -- $08691
          34450 => x"80", -- $08692
          34451 => x"80", -- $08693
          34452 => x"80", -- $08694
          34453 => x"80", -- $08695
          34454 => x"80", -- $08696
          34455 => x"80", -- $08697
          34456 => x"80", -- $08698
          34457 => x"80", -- $08699
          34458 => x"80", -- $0869a
          34459 => x"80", -- $0869b
          34460 => x"80", -- $0869c
          34461 => x"80", -- $0869d
          34462 => x"80", -- $0869e
          34463 => x"80", -- $0869f
          34464 => x"80", -- $086a0
          34465 => x"80", -- $086a1
          34466 => x"80", -- $086a2
          34467 => x"80", -- $086a3
          34468 => x"80", -- $086a4
          34469 => x"80", -- $086a5
          34470 => x"80", -- $086a6
          34471 => x"80", -- $086a7
          34472 => x"80", -- $086a8
          34473 => x"80", -- $086a9
          34474 => x"80", -- $086aa
          34475 => x"80", -- $086ab
          34476 => x"80", -- $086ac
          34477 => x"80", -- $086ad
          34478 => x"80", -- $086ae
          34479 => x"80", -- $086af
          34480 => x"80", -- $086b0
          34481 => x"80", -- $086b1
          34482 => x"80", -- $086b2
          34483 => x"80", -- $086b3
          34484 => x"80", -- $086b4
          34485 => x"80", -- $086b5
          34486 => x"80", -- $086b6
          34487 => x"80", -- $086b7
          34488 => x"80", -- $086b8
          34489 => x"80", -- $086b9
          34490 => x"80", -- $086ba
          34491 => x"80", -- $086bb
          34492 => x"80", -- $086bc
          34493 => x"80", -- $086bd
          34494 => x"80", -- $086be
          34495 => x"80", -- $086bf
          34496 => x"80", -- $086c0
          34497 => x"80", -- $086c1
          34498 => x"80", -- $086c2
          34499 => x"81", -- $086c3
          34500 => x"81", -- $086c4
          34501 => x"81", -- $086c5
          34502 => x"81", -- $086c6
          34503 => x"81", -- $086c7
          34504 => x"81", -- $086c8
          34505 => x"81", -- $086c9
          34506 => x"81", -- $086ca
          34507 => x"80", -- $086cb
          34508 => x"80", -- $086cc
          34509 => x"80", -- $086cd
          34510 => x"80", -- $086ce
          34511 => x"80", -- $086cf
          34512 => x"80", -- $086d0
          34513 => x"80", -- $086d1
          34514 => x"80", -- $086d2
          34515 => x"80", -- $086d3
          34516 => x"80", -- $086d4
          34517 => x"80", -- $086d5
          34518 => x"80", -- $086d6
          34519 => x"80", -- $086d7
          34520 => x"80", -- $086d8
          34521 => x"80", -- $086d9
          34522 => x"80", -- $086da
          34523 => x"80", -- $086db
          34524 => x"81", -- $086dc
          34525 => x"81", -- $086dd
          34526 => x"81", -- $086de
          34527 => x"81", -- $086df
          34528 => x"81", -- $086e0
          34529 => x"81", -- $086e1
          34530 => x"81", -- $086e2
          34531 => x"81", -- $086e3
          34532 => x"81", -- $086e4
          34533 => x"81", -- $086e5
          34534 => x"81", -- $086e6
          34535 => x"81", -- $086e7
          34536 => x"81", -- $086e8
          34537 => x"81", -- $086e9
          34538 => x"81", -- $086ea
          34539 => x"81", -- $086eb
          34540 => x"81", -- $086ec
          34541 => x"81", -- $086ed
          34542 => x"81", -- $086ee
          34543 => x"81", -- $086ef
          34544 => x"81", -- $086f0
          34545 => x"81", -- $086f1
          34546 => x"81", -- $086f2
          34547 => x"81", -- $086f3
          34548 => x"80", -- $086f4
          34549 => x"80", -- $086f5
          34550 => x"80", -- $086f6
          34551 => x"81", -- $086f7
          34552 => x"81", -- $086f8
          34553 => x"81", -- $086f9
          34554 => x"81", -- $086fa
          34555 => x"81", -- $086fb
          34556 => x"81", -- $086fc
          34557 => x"81", -- $086fd
          34558 => x"81", -- $086fe
          34559 => x"81", -- $086ff
          34560 => x"81", -- $08700
          34561 => x"81", -- $08701
          34562 => x"81", -- $08702
          34563 => x"82", -- $08703
          34564 => x"82", -- $08704
          34565 => x"82", -- $08705
          34566 => x"82", -- $08706
          34567 => x"82", -- $08707
          34568 => x"82", -- $08708
          34569 => x"82", -- $08709
          34570 => x"82", -- $0870a
          34571 => x"82", -- $0870b
          34572 => x"82", -- $0870c
          34573 => x"82", -- $0870d
          34574 => x"82", -- $0870e
          34575 => x"81", -- $0870f
          34576 => x"81", -- $08710
          34577 => x"81", -- $08711
          34578 => x"81", -- $08712
          34579 => x"81", -- $08713
          34580 => x"81", -- $08714
          34581 => x"81", -- $08715
          34582 => x"81", -- $08716
          34583 => x"81", -- $08717
          34584 => x"81", -- $08718
          34585 => x"81", -- $08719
          34586 => x"81", -- $0871a
          34587 => x"81", -- $0871b
          34588 => x"81", -- $0871c
          34589 => x"81", -- $0871d
          34590 => x"81", -- $0871e
          34591 => x"81", -- $0871f
          34592 => x"82", -- $08720
          34593 => x"82", -- $08721
          34594 => x"82", -- $08722
          34595 => x"82", -- $08723
          34596 => x"82", -- $08724
          34597 => x"82", -- $08725
          34598 => x"82", -- $08726
          34599 => x"82", -- $08727
          34600 => x"82", -- $08728
          34601 => x"82", -- $08729
          34602 => x"82", -- $0872a
          34603 => x"82", -- $0872b
          34604 => x"82", -- $0872c
          34605 => x"82", -- $0872d
          34606 => x"82", -- $0872e
          34607 => x"82", -- $0872f
          34608 => x"82", -- $08730
          34609 => x"82", -- $08731
          34610 => x"81", -- $08732
          34611 => x"81", -- $08733
          34612 => x"81", -- $08734
          34613 => x"81", -- $08735
          34614 => x"81", -- $08736
          34615 => x"81", -- $08737
          34616 => x"81", -- $08738
          34617 => x"81", -- $08739
          34618 => x"81", -- $0873a
          34619 => x"81", -- $0873b
          34620 => x"81", -- $0873c
          34621 => x"81", -- $0873d
          34622 => x"81", -- $0873e
          34623 => x"81", -- $0873f
          34624 => x"81", -- $08740
          34625 => x"82", -- $08741
          34626 => x"82", -- $08742
          34627 => x"82", -- $08743
          34628 => x"82", -- $08744
          34629 => x"82", -- $08745
          34630 => x"82", -- $08746
          34631 => x"82", -- $08747
          34632 => x"82", -- $08748
          34633 => x"82", -- $08749
          34634 => x"82", -- $0874a
          34635 => x"82", -- $0874b
          34636 => x"82", -- $0874c
          34637 => x"82", -- $0874d
          34638 => x"82", -- $0874e
          34639 => x"82", -- $0874f
          34640 => x"82", -- $08750
          34641 => x"81", -- $08751
          34642 => x"81", -- $08752
          34643 => x"81", -- $08753
          34644 => x"81", -- $08754
          34645 => x"81", -- $08755
          34646 => x"81", -- $08756
          34647 => x"81", -- $08757
          34648 => x"81", -- $08758
          34649 => x"81", -- $08759
          34650 => x"81", -- $0875a
          34651 => x"81", -- $0875b
          34652 => x"81", -- $0875c
          34653 => x"81", -- $0875d
          34654 => x"81", -- $0875e
          34655 => x"81", -- $0875f
          34656 => x"81", -- $08760
          34657 => x"81", -- $08761
          34658 => x"81", -- $08762
          34659 => x"81", -- $08763
          34660 => x"81", -- $08764
          34661 => x"81", -- $08765
          34662 => x"81", -- $08766
          34663 => x"81", -- $08767
          34664 => x"81", -- $08768
          34665 => x"81", -- $08769
          34666 => x"81", -- $0876a
          34667 => x"81", -- $0876b
          34668 => x"81", -- $0876c
          34669 => x"81", -- $0876d
          34670 => x"81", -- $0876e
          34671 => x"81", -- $0876f
          34672 => x"81", -- $08770
          34673 => x"81", -- $08771
          34674 => x"81", -- $08772
          34675 => x"81", -- $08773
          34676 => x"81", -- $08774
          34677 => x"81", -- $08775
          34678 => x"80", -- $08776
          34679 => x"80", -- $08777
          34680 => x"80", -- $08778
          34681 => x"80", -- $08779
          34682 => x"80", -- $0877a
          34683 => x"80", -- $0877b
          34684 => x"80", -- $0877c
          34685 => x"80", -- $0877d
          34686 => x"80", -- $0877e
          34687 => x"80", -- $0877f
          34688 => x"80", -- $08780
          34689 => x"80", -- $08781
          34690 => x"80", -- $08782
          34691 => x"80", -- $08783
          34692 => x"80", -- $08784
          34693 => x"80", -- $08785
          34694 => x"80", -- $08786
          34695 => x"81", -- $08787
          34696 => x"81", -- $08788
          34697 => x"81", -- $08789
          34698 => x"81", -- $0878a
          34699 => x"81", -- $0878b
          34700 => x"81", -- $0878c
          34701 => x"81", -- $0878d
          34702 => x"81", -- $0878e
          34703 => x"81", -- $0878f
          34704 => x"81", -- $08790
          34705 => x"81", -- $08791
          34706 => x"81", -- $08792
          34707 => x"81", -- $08793
          34708 => x"80", -- $08794
          34709 => x"80", -- $08795
          34710 => x"80", -- $08796
          34711 => x"80", -- $08797
          34712 => x"80", -- $08798
          34713 => x"80", -- $08799
          34714 => x"80", -- $0879a
          34715 => x"80", -- $0879b
          34716 => x"80", -- $0879c
          34717 => x"80", -- $0879d
          34718 => x"80", -- $0879e
          34719 => x"80", -- $0879f
          34720 => x"80", -- $087a0
          34721 => x"80", -- $087a1
          34722 => x"80", -- $087a2
          34723 => x"80", -- $087a3
          34724 => x"80", -- $087a4
          34725 => x"80", -- $087a5
          34726 => x"80", -- $087a6
          34727 => x"80", -- $087a7
          34728 => x"80", -- $087a8
          34729 => x"80", -- $087a9
          34730 => x"80", -- $087aa
          34731 => x"80", -- $087ab
          34732 => x"80", -- $087ac
          34733 => x"80", -- $087ad
          34734 => x"80", -- $087ae
          34735 => x"80", -- $087af
          34736 => x"81", -- $087b0
          34737 => x"81", -- $087b1
          34738 => x"80", -- $087b2
          34739 => x"80", -- $087b3
          34740 => x"80", -- $087b4
          34741 => x"80", -- $087b5
          34742 => x"80", -- $087b6
          34743 => x"80", -- $087b7
          34744 => x"80", -- $087b8
          34745 => x"80", -- $087b9
          34746 => x"80", -- $087ba
          34747 => x"80", -- $087bb
          34748 => x"80", -- $087bc
          34749 => x"80", -- $087bd
          34750 => x"80", -- $087be
          34751 => x"80", -- $087bf
          34752 => x"80", -- $087c0
          34753 => x"80", -- $087c1
          34754 => x"80", -- $087c2
          34755 => x"80", -- $087c3
          34756 => x"80", -- $087c4
          34757 => x"80", -- $087c5
          34758 => x"80", -- $087c6
          34759 => x"80", -- $087c7
          34760 => x"80", -- $087c8
          34761 => x"80", -- $087c9
          34762 => x"80", -- $087ca
          34763 => x"80", -- $087cb
          34764 => x"80", -- $087cc
          34765 => x"80", -- $087cd
          34766 => x"80", -- $087ce
          34767 => x"80", -- $087cf
          34768 => x"81", -- $087d0
          34769 => x"81", -- $087d1
          34770 => x"81", -- $087d2
          34771 => x"81", -- $087d3
          34772 => x"81", -- $087d4
          34773 => x"81", -- $087d5
          34774 => x"81", -- $087d6
          34775 => x"80", -- $087d7
          34776 => x"80", -- $087d8
          34777 => x"80", -- $087d9
          34778 => x"80", -- $087da
          34779 => x"80", -- $087db
          34780 => x"80", -- $087dc
          34781 => x"80", -- $087dd
          34782 => x"80", -- $087de
          34783 => x"80", -- $087df
          34784 => x"80", -- $087e0
          34785 => x"80", -- $087e1
          34786 => x"80", -- $087e2
          34787 => x"80", -- $087e3
          34788 => x"80", -- $087e4
          34789 => x"80", -- $087e5
          34790 => x"80", -- $087e6
          34791 => x"80", -- $087e7
          34792 => x"80", -- $087e8
          34793 => x"80", -- $087e9
          34794 => x"80", -- $087ea
          34795 => x"80", -- $087eb
          34796 => x"80", -- $087ec
          34797 => x"80", -- $087ed
          34798 => x"80", -- $087ee
          34799 => x"80", -- $087ef
          34800 => x"80", -- $087f0
          34801 => x"80", -- $087f1
          34802 => x"80", -- $087f2
          34803 => x"80", -- $087f3
          34804 => x"80", -- $087f4
          34805 => x"80", -- $087f5
          34806 => x"80", -- $087f6
          34807 => x"80", -- $087f7
          34808 => x"80", -- $087f8
          34809 => x"80", -- $087f9
          34810 => x"80", -- $087fa
          34811 => x"80", -- $087fb
          34812 => x"80", -- $087fc
          34813 => x"80", -- $087fd
          34814 => x"80", -- $087fe
          34815 => x"80", -- $087ff
          34816 => x"80", -- $08800
          34817 => x"80", -- $08801
          34818 => x"80", -- $08802
          34819 => x"80", -- $08803
          34820 => x"80", -- $08804
          34821 => x"80", -- $08805
          34822 => x"80", -- $08806
          34823 => x"80", -- $08807
          34824 => x"80", -- $08808
          34825 => x"80", -- $08809
          34826 => x"80", -- $0880a
          34827 => x"80", -- $0880b
          34828 => x"80", -- $0880c
          34829 => x"80", -- $0880d
          34830 => x"80", -- $0880e
          34831 => x"80", -- $0880f
          34832 => x"80", -- $08810
          34833 => x"80", -- $08811
          34834 => x"80", -- $08812
          34835 => x"80", -- $08813
          34836 => x"80", -- $08814
          34837 => x"80", -- $08815
          34838 => x"80", -- $08816
          34839 => x"80", -- $08817
          34840 => x"80", -- $08818
          34841 => x"80", -- $08819
          34842 => x"80", -- $0881a
          34843 => x"80", -- $0881b
          34844 => x"80", -- $0881c
          34845 => x"80", -- $0881d
          34846 => x"80", -- $0881e
          34847 => x"80", -- $0881f
          34848 => x"7f", -- $08820
          34849 => x"7f", -- $08821
          34850 => x"7f", -- $08822
          34851 => x"7f", -- $08823
          34852 => x"7f", -- $08824
          34853 => x"7f", -- $08825
          34854 => x"7f", -- $08826
          34855 => x"7f", -- $08827
          34856 => x"7f", -- $08828
          34857 => x"7f", -- $08829
          34858 => x"7f", -- $0882a
          34859 => x"7f", -- $0882b
          34860 => x"7f", -- $0882c
          34861 => x"7f", -- $0882d
          34862 => x"80", -- $0882e
          34863 => x"80", -- $0882f
          34864 => x"80", -- $08830
          34865 => x"80", -- $08831
          34866 => x"80", -- $08832
          34867 => x"80", -- $08833
          34868 => x"80", -- $08834
          34869 => x"80", -- $08835
          34870 => x"80", -- $08836
          34871 => x"80", -- $08837
          34872 => x"80", -- $08838
          34873 => x"80", -- $08839
          34874 => x"80", -- $0883a
          34875 => x"7f", -- $0883b
          34876 => x"7f", -- $0883c
          34877 => x"7f", -- $0883d
          34878 => x"7f", -- $0883e
          34879 => x"7f", -- $0883f
          34880 => x"7f", -- $08840
          34881 => x"7f", -- $08841
          34882 => x"7f", -- $08842
          34883 => x"7f", -- $08843
          34884 => x"7f", -- $08844
          34885 => x"7f", -- $08845
          34886 => x"7f", -- $08846
          34887 => x"7f", -- $08847
          34888 => x"7f", -- $08848
          34889 => x"7f", -- $08849
          34890 => x"7f", -- $0884a
          34891 => x"7f", -- $0884b
          34892 => x"7f", -- $0884c
          34893 => x"7f", -- $0884d
          34894 => x"7f", -- $0884e
          34895 => x"7f", -- $0884f
          34896 => x"7f", -- $08850
          34897 => x"7f", -- $08851
          34898 => x"7f", -- $08852
          34899 => x"7f", -- $08853
          34900 => x"7f", -- $08854
          34901 => x"7f", -- $08855
          34902 => x"7f", -- $08856
          34903 => x"7f", -- $08857
          34904 => x"7f", -- $08858
          34905 => x"7f", -- $08859
          34906 => x"7f", -- $0885a
          34907 => x"7f", -- $0885b
          34908 => x"7f", -- $0885c
          34909 => x"7f", -- $0885d
          34910 => x"7f", -- $0885e
          34911 => x"7f", -- $0885f
          34912 => x"7f", -- $08860
          34913 => x"7f", -- $08861
          34914 => x"7f", -- $08862
          34915 => x"7f", -- $08863
          34916 => x"7f", -- $08864
          34917 => x"7f", -- $08865
          34918 => x"7f", -- $08866
          34919 => x"7f", -- $08867
          34920 => x"7f", -- $08868
          34921 => x"7f", -- $08869
          34922 => x"7f", -- $0886a
          34923 => x"7f", -- $0886b
          34924 => x"7f", -- $0886c
          34925 => x"7f", -- $0886d
          34926 => x"7f", -- $0886e
          34927 => x"7f", -- $0886f
          34928 => x"7f", -- $08870
          34929 => x"7f", -- $08871
          34930 => x"7f", -- $08872
          34931 => x"7f", -- $08873
          34932 => x"7f", -- $08874
          34933 => x"7f", -- $08875
          34934 => x"7f", -- $08876
          34935 => x"7f", -- $08877
          34936 => x"7f", -- $08878
          34937 => x"7f", -- $08879
          34938 => x"7f", -- $0887a
          34939 => x"7f", -- $0887b
          34940 => x"7f", -- $0887c
          34941 => x"7f", -- $0887d
          34942 => x"7f", -- $0887e
          34943 => x"7f", -- $0887f
          34944 => x"7f", -- $08880
          34945 => x"7f", -- $08881
          34946 => x"7f", -- $08882
          34947 => x"7f", -- $08883
          34948 => x"7f", -- $08884
          34949 => x"7f", -- $08885
          34950 => x"7e", -- $08886
          34951 => x"7e", -- $08887
          34952 => x"7e", -- $08888
          34953 => x"7f", -- $08889
          34954 => x"7f", -- $0888a
          34955 => x"7f", -- $0888b
          34956 => x"7f", -- $0888c
          34957 => x"7f", -- $0888d
          34958 => x"7f", -- $0888e
          34959 => x"7f", -- $0888f
          34960 => x"7f", -- $08890
          34961 => x"7f", -- $08891
          34962 => x"7f", -- $08892
          34963 => x"7f", -- $08893
          34964 => x"7f", -- $08894
          34965 => x"7f", -- $08895
          34966 => x"7f", -- $08896
          34967 => x"7f", -- $08897
          34968 => x"7f", -- $08898
          34969 => x"7f", -- $08899
          34970 => x"7f", -- $0889a
          34971 => x"7f", -- $0889b
          34972 => x"7f", -- $0889c
          34973 => x"7f", -- $0889d
          34974 => x"7f", -- $0889e
          34975 => x"7f", -- $0889f
          34976 => x"7f", -- $088a0
          34977 => x"7f", -- $088a1
          34978 => x"7f", -- $088a2
          34979 => x"7f", -- $088a3
          34980 => x"7f", -- $088a4
          34981 => x"7f", -- $088a5
          34982 => x"7f", -- $088a6
          34983 => x"7f", -- $088a7
          34984 => x"7f", -- $088a8
          34985 => x"7f", -- $088a9
          34986 => x"7f", -- $088aa
          34987 => x"7f", -- $088ab
          34988 => x"7f", -- $088ac
          34989 => x"7f", -- $088ad
          34990 => x"7f", -- $088ae
          34991 => x"7f", -- $088af
          34992 => x"7f", -- $088b0
          34993 => x"7f", -- $088b1
          34994 => x"7f", -- $088b2
          34995 => x"7f", -- $088b3
          34996 => x"80", -- $088b4
          34997 => x"80", -- $088b5
          34998 => x"80", -- $088b6
          34999 => x"80", -- $088b7
          35000 => x"80", -- $088b8
          35001 => x"80", -- $088b9
          35002 => x"7f", -- $088ba
          35003 => x"7f", -- $088bb
          35004 => x"7f", -- $088bc
          35005 => x"7f", -- $088bd
          35006 => x"7f", -- $088be
          35007 => x"7f", -- $088bf
          35008 => x"7f", -- $088c0
          35009 => x"7f", -- $088c1
          35010 => x"7f", -- $088c2
          35011 => x"7f", -- $088c3
          35012 => x"7f", -- $088c4
          35013 => x"7f", -- $088c5
          35014 => x"7f", -- $088c6
          35015 => x"7f", -- $088c7
          35016 => x"7f", -- $088c8
          35017 => x"7f", -- $088c9
          35018 => x"7f", -- $088ca
          35019 => x"7f", -- $088cb
          35020 => x"7f", -- $088cc
          35021 => x"7f", -- $088cd
          35022 => x"7f", -- $088ce
          35023 => x"80", -- $088cf
          35024 => x"80", -- $088d0
          35025 => x"80", -- $088d1
          35026 => x"80", -- $088d2
          35027 => x"80", -- $088d3
          35028 => x"80", -- $088d4
          35029 => x"80", -- $088d5
          35030 => x"80", -- $088d6
          35031 => x"80", -- $088d7
          35032 => x"80", -- $088d8
          35033 => x"80", -- $088d9
          35034 => x"80", -- $088da
          35035 => x"80", -- $088db
          35036 => x"7f", -- $088dc
          35037 => x"7f", -- $088dd
          35038 => x"7f", -- $088de
          35039 => x"7f", -- $088df
          35040 => x"7f", -- $088e0
          35041 => x"7f", -- $088e1
          35042 => x"7f", -- $088e2
          35043 => x"7f", -- $088e3
          35044 => x"7f", -- $088e4
          35045 => x"7f", -- $088e5
          35046 => x"7f", -- $088e6
          35047 => x"7f", -- $088e7
          35048 => x"7f", -- $088e8
          35049 => x"7f", -- $088e9
          35050 => x"7f", -- $088ea
          35051 => x"7f", -- $088eb
          35052 => x"7f", -- $088ec
          35053 => x"7f", -- $088ed
          35054 => x"7f", -- $088ee
          35055 => x"7f", -- $088ef
          35056 => x"7f", -- $088f0
          35057 => x"80", -- $088f1
          35058 => x"80", -- $088f2
          35059 => x"80", -- $088f3
          35060 => x"80", -- $088f4
          35061 => x"80", -- $088f5
          35062 => x"80", -- $088f6
          35063 => x"80", -- $088f7
          35064 => x"80", -- $088f8
          35065 => x"80", -- $088f9
          35066 => x"80", -- $088fa
          35067 => x"7f", -- $088fb
          35068 => x"7f", -- $088fc
          35069 => x"7f", -- $088fd
          35070 => x"7f", -- $088fe
          35071 => x"7f", -- $088ff
          35072 => x"7f", -- $08900
          35073 => x"7f", -- $08901
          35074 => x"7f", -- $08902
          35075 => x"7f", -- $08903
          35076 => x"7f", -- $08904
          35077 => x"7f", -- $08905
          35078 => x"7f", -- $08906
          35079 => x"7f", -- $08907
          35080 => x"7f", -- $08908
          35081 => x"7f", -- $08909
          35082 => x"7f", -- $0890a
          35083 => x"7f", -- $0890b
          35084 => x"7f", -- $0890c
          35085 => x"7f", -- $0890d
          35086 => x"80", -- $0890e
          35087 => x"80", -- $0890f
          35088 => x"80", -- $08910
          35089 => x"80", -- $08911
          35090 => x"80", -- $08912
          35091 => x"80", -- $08913
          35092 => x"80", -- $08914
          35093 => x"80", -- $08915
          35094 => x"80", -- $08916
          35095 => x"80", -- $08917
          35096 => x"80", -- $08918
          35097 => x"80", -- $08919
          35098 => x"80", -- $0891a
          35099 => x"7f", -- $0891b
          35100 => x"7f", -- $0891c
          35101 => x"7f", -- $0891d
          35102 => x"7f", -- $0891e
          35103 => x"7f", -- $0891f
          35104 => x"7f", -- $08920
          35105 => x"7f", -- $08921
          35106 => x"7f", -- $08922
          35107 => x"7f", -- $08923
          35108 => x"7f", -- $08924
          35109 => x"7f", -- $08925
          35110 => x"7f", -- $08926
          35111 => x"7f", -- $08927
          35112 => x"7f", -- $08928
          35113 => x"7f", -- $08929
          35114 => x"80", -- $0892a
          35115 => x"80", -- $0892b
          35116 => x"80", -- $0892c
          35117 => x"80", -- $0892d
          35118 => x"80", -- $0892e
          35119 => x"80", -- $0892f
          35120 => x"80", -- $08930
          35121 => x"80", -- $08931
          35122 => x"80", -- $08932
          35123 => x"80", -- $08933
          35124 => x"80", -- $08934
          35125 => x"80", -- $08935
          35126 => x"80", -- $08936
          35127 => x"80", -- $08937
          35128 => x"80", -- $08938
          35129 => x"80", -- $08939
          35130 => x"80", -- $0893a
          35131 => x"80", -- $0893b
          35132 => x"80", -- $0893c
          35133 => x"80", -- $0893d
          35134 => x"80", -- $0893e
          35135 => x"80", -- $0893f
          35136 => x"80", -- $08940
          35137 => x"80", -- $08941
          35138 => x"80", -- $08942
          35139 => x"7f", -- $08943
          35140 => x"80", -- $08944
          35141 => x"80", -- $08945
          35142 => x"80", -- $08946
          35143 => x"80", -- $08947
          35144 => x"80", -- $08948
          35145 => x"80", -- $08949
          35146 => x"80", -- $0894a
          35147 => x"80", -- $0894b
          35148 => x"80", -- $0894c
          35149 => x"80", -- $0894d
          35150 => x"80", -- $0894e
          35151 => x"80", -- $0894f
          35152 => x"80", -- $08950
          35153 => x"80", -- $08951
          35154 => x"80", -- $08952
          35155 => x"80", -- $08953
          35156 => x"80", -- $08954
          35157 => x"80", -- $08955
          35158 => x"80", -- $08956
          35159 => x"80", -- $08957
          35160 => x"80", -- $08958
          35161 => x"80", -- $08959
          35162 => x"80", -- $0895a
          35163 => x"80", -- $0895b
          35164 => x"80", -- $0895c
          35165 => x"80", -- $0895d
          35166 => x"80", -- $0895e
          35167 => x"80", -- $0895f
          35168 => x"80", -- $08960
          35169 => x"80", -- $08961
          35170 => x"80", -- $08962
          35171 => x"80", -- $08963
          35172 => x"80", -- $08964
          35173 => x"80", -- $08965
          35174 => x"80", -- $08966
          35175 => x"80", -- $08967
          35176 => x"80", -- $08968
          35177 => x"80", -- $08969
          35178 => x"80", -- $0896a
          35179 => x"80", -- $0896b
          35180 => x"80", -- $0896c
          35181 => x"80", -- $0896d
          35182 => x"80", -- $0896e
          35183 => x"80", -- $0896f
          35184 => x"80", -- $08970
          35185 => x"80", -- $08971
          35186 => x"80", -- $08972
          35187 => x"80", -- $08973
          35188 => x"80", -- $08974
          35189 => x"80", -- $08975
          35190 => x"80", -- $08976
          35191 => x"80", -- $08977
          35192 => x"80", -- $08978
          35193 => x"80", -- $08979
          35194 => x"80", -- $0897a
          35195 => x"80", -- $0897b
          35196 => x"80", -- $0897c
          35197 => x"80", -- $0897d
          35198 => x"80", -- $0897e
          35199 => x"80", -- $0897f
          35200 => x"80", -- $08980
          35201 => x"80", -- $08981
          35202 => x"80", -- $08982
          35203 => x"80", -- $08983
          35204 => x"80", -- $08984
          35205 => x"80", -- $08985
          35206 => x"80", -- $08986
          35207 => x"80", -- $08987
          35208 => x"80", -- $08988
          35209 => x"80", -- $08989
          35210 => x"80", -- $0898a
          35211 => x"80", -- $0898b
          35212 => x"80", -- $0898c
          35213 => x"80", -- $0898d
          35214 => x"80", -- $0898e
          35215 => x"80", -- $0898f
          35216 => x"81", -- $08990
          35217 => x"81", -- $08991
          35218 => x"81", -- $08992
          35219 => x"81", -- $08993
          35220 => x"81", -- $08994
          35221 => x"81", -- $08995
          35222 => x"80", -- $08996
          35223 => x"80", -- $08997
          35224 => x"80", -- $08998
          35225 => x"80", -- $08999
          35226 => x"80", -- $0899a
          35227 => x"80", -- $0899b
          35228 => x"80", -- $0899c
          35229 => x"80", -- $0899d
          35230 => x"80", -- $0899e
          35231 => x"80", -- $0899f
          35232 => x"80", -- $089a0
          35233 => x"80", -- $089a1
          35234 => x"80", -- $089a2
          35235 => x"80", -- $089a3
          35236 => x"80", -- $089a4
          35237 => x"80", -- $089a5
          35238 => x"80", -- $089a6
          35239 => x"80", -- $089a7
          35240 => x"80", -- $089a8
          35241 => x"80", -- $089a9
          35242 => x"80", -- $089aa
          35243 => x"80", -- $089ab
          35244 => x"80", -- $089ac
          35245 => x"80", -- $089ad
          35246 => x"80", -- $089ae
          35247 => x"81", -- $089af
          35248 => x"81", -- $089b0
          35249 => x"81", -- $089b1
          35250 => x"81", -- $089b2
          35251 => x"81", -- $089b3
          35252 => x"81", -- $089b4
          35253 => x"81", -- $089b5
          35254 => x"80", -- $089b6
          35255 => x"80", -- $089b7
          35256 => x"80", -- $089b8
          35257 => x"80", -- $089b9
          35258 => x"80", -- $089ba
          35259 => x"80", -- $089bb
          35260 => x"80", -- $089bc
          35261 => x"80", -- $089bd
          35262 => x"80", -- $089be
          35263 => x"80", -- $089bf
          35264 => x"80", -- $089c0
          35265 => x"80", -- $089c1
          35266 => x"80", -- $089c2
          35267 => x"80", -- $089c3
          35268 => x"80", -- $089c4
          35269 => x"80", -- $089c5
          35270 => x"80", -- $089c6
          35271 => x"81", -- $089c7
          35272 => x"81", -- $089c8
          35273 => x"81", -- $089c9
          35274 => x"81", -- $089ca
          35275 => x"81", -- $089cb
          35276 => x"81", -- $089cc
          35277 => x"81", -- $089cd
          35278 => x"81", -- $089ce
          35279 => x"81", -- $089cf
          35280 => x"81", -- $089d0
          35281 => x"81", -- $089d1
          35282 => x"81", -- $089d2
          35283 => x"81", -- $089d3
          35284 => x"81", -- $089d4
          35285 => x"81", -- $089d5
          35286 => x"81", -- $089d6
          35287 => x"81", -- $089d7
          35288 => x"81", -- $089d8
          35289 => x"81", -- $089d9
          35290 => x"80", -- $089da
          35291 => x"80", -- $089db
          35292 => x"80", -- $089dc
          35293 => x"80", -- $089dd
          35294 => x"80", -- $089de
          35295 => x"80", -- $089df
          35296 => x"80", -- $089e0
          35297 => x"80", -- $089e1
          35298 => x"80", -- $089e2
          35299 => x"80", -- $089e3
          35300 => x"80", -- $089e4
          35301 => x"80", -- $089e5
          35302 => x"81", -- $089e6
          35303 => x"81", -- $089e7
          35304 => x"81", -- $089e8
          35305 => x"81", -- $089e9
          35306 => x"81", -- $089ea
          35307 => x"81", -- $089eb
          35308 => x"81", -- $089ec
          35309 => x"81", -- $089ed
          35310 => x"81", -- $089ee
          35311 => x"81", -- $089ef
          35312 => x"81", -- $089f0
          35313 => x"81", -- $089f1
          35314 => x"81", -- $089f2
          35315 => x"80", -- $089f3
          35316 => x"80", -- $089f4
          35317 => x"80", -- $089f5
          35318 => x"80", -- $089f6
          35319 => x"80", -- $089f7
          35320 => x"80", -- $089f8
          35321 => x"80", -- $089f9
          35322 => x"80", -- $089fa
          35323 => x"80", -- $089fb
          35324 => x"80", -- $089fc
          35325 => x"80", -- $089fd
          35326 => x"80", -- $089fe
          35327 => x"80", -- $089ff
          35328 => x"80", -- $08a00
          35329 => x"80", -- $08a01
          35330 => x"80", -- $08a02
          35331 => x"80", -- $08a03
          35332 => x"80", -- $08a04
          35333 => x"80", -- $08a05
          35334 => x"80", -- $08a06
          35335 => x"80", -- $08a07
          35336 => x"80", -- $08a08
          35337 => x"81", -- $08a09
          35338 => x"81", -- $08a0a
          35339 => x"80", -- $08a0b
          35340 => x"80", -- $08a0c
          35341 => x"80", -- $08a0d
          35342 => x"80", -- $08a0e
          35343 => x"80", -- $08a0f
          35344 => x"80", -- $08a10
          35345 => x"80", -- $08a11
          35346 => x"80", -- $08a12
          35347 => x"80", -- $08a13
          35348 => x"80", -- $08a14
          35349 => x"80", -- $08a15
          35350 => x"80", -- $08a16
          35351 => x"80", -- $08a17
          35352 => x"80", -- $08a18
          35353 => x"80", -- $08a19
          35354 => x"80", -- $08a1a
          35355 => x"80", -- $08a1b
          35356 => x"80", -- $08a1c
          35357 => x"80", -- $08a1d
          35358 => x"80", -- $08a1e
          35359 => x"80", -- $08a1f
          35360 => x"80", -- $08a20
          35361 => x"80", -- $08a21
          35362 => x"80", -- $08a22
          35363 => x"80", -- $08a23
          35364 => x"80", -- $08a24
          35365 => x"80", -- $08a25
          35366 => x"80", -- $08a26
          35367 => x"80", -- $08a27
          35368 => x"80", -- $08a28
          35369 => x"80", -- $08a29
          35370 => x"80", -- $08a2a
          35371 => x"80", -- $08a2b
          35372 => x"80", -- $08a2c
          35373 => x"80", -- $08a2d
          35374 => x"80", -- $08a2e
          35375 => x"81", -- $08a2f
          35376 => x"81", -- $08a30
          35377 => x"81", -- $08a31
          35378 => x"81", -- $08a32
          35379 => x"81", -- $08a33
          35380 => x"81", -- $08a34
          35381 => x"81", -- $08a35
          35382 => x"81", -- $08a36
          35383 => x"81", -- $08a37
          35384 => x"81", -- $08a38
          35385 => x"81", -- $08a39
          35386 => x"80", -- $08a3a
          35387 => x"81", -- $08a3b
          35388 => x"81", -- $08a3c
          35389 => x"81", -- $08a3d
          35390 => x"81", -- $08a3e
          35391 => x"81", -- $08a3f
          35392 => x"81", -- $08a40
          35393 => x"81", -- $08a41
          35394 => x"81", -- $08a42
          35395 => x"81", -- $08a43
          35396 => x"81", -- $08a44
          35397 => x"81", -- $08a45
          35398 => x"81", -- $08a46
          35399 => x"81", -- $08a47
          35400 => x"81", -- $08a48
          35401 => x"81", -- $08a49
          35402 => x"81", -- $08a4a
          35403 => x"81", -- $08a4b
          35404 => x"81", -- $08a4c
          35405 => x"81", -- $08a4d
          35406 => x"81", -- $08a4e
          35407 => x"81", -- $08a4f
          35408 => x"81", -- $08a50
          35409 => x"81", -- $08a51
          35410 => x"81", -- $08a52
          35411 => x"81", -- $08a53
          35412 => x"81", -- $08a54
          35413 => x"81", -- $08a55
          35414 => x"81", -- $08a56
          35415 => x"81", -- $08a57
          35416 => x"81", -- $08a58
          35417 => x"81", -- $08a59
          35418 => x"81", -- $08a5a
          35419 => x"81", -- $08a5b
          35420 => x"81", -- $08a5c
          35421 => x"81", -- $08a5d
          35422 => x"81", -- $08a5e
          35423 => x"81", -- $08a5f
          35424 => x"81", -- $08a60
          35425 => x"81", -- $08a61
          35426 => x"81", -- $08a62
          35427 => x"81", -- $08a63
          35428 => x"81", -- $08a64
          35429 => x"81", -- $08a65
          35430 => x"81", -- $08a66
          35431 => x"81", -- $08a67
          35432 => x"81", -- $08a68
          35433 => x"81", -- $08a69
          35434 => x"81", -- $08a6a
          35435 => x"81", -- $08a6b
          35436 => x"81", -- $08a6c
          35437 => x"81", -- $08a6d
          35438 => x"81", -- $08a6e
          35439 => x"81", -- $08a6f
          35440 => x"81", -- $08a70
          35441 => x"81", -- $08a71
          35442 => x"81", -- $08a72
          35443 => x"81", -- $08a73
          35444 => x"81", -- $08a74
          35445 => x"81", -- $08a75
          35446 => x"81", -- $08a76
          35447 => x"81", -- $08a77
          35448 => x"81", -- $08a78
          35449 => x"81", -- $08a79
          35450 => x"81", -- $08a7a
          35451 => x"81", -- $08a7b
          35452 => x"81", -- $08a7c
          35453 => x"81", -- $08a7d
          35454 => x"81", -- $08a7e
          35455 => x"81", -- $08a7f
          35456 => x"81", -- $08a80
          35457 => x"81", -- $08a81
          35458 => x"80", -- $08a82
          35459 => x"80", -- $08a83
          35460 => x"80", -- $08a84
          35461 => x"80", -- $08a85
          35462 => x"80", -- $08a86
          35463 => x"80", -- $08a87
          35464 => x"80", -- $08a88
          35465 => x"80", -- $08a89
          35466 => x"80", -- $08a8a
          35467 => x"80", -- $08a8b
          35468 => x"81", -- $08a8c
          35469 => x"81", -- $08a8d
          35470 => x"80", -- $08a8e
          35471 => x"80", -- $08a8f
          35472 => x"80", -- $08a90
          35473 => x"80", -- $08a91
          35474 => x"80", -- $08a92
          35475 => x"80", -- $08a93
          35476 => x"80", -- $08a94
          35477 => x"80", -- $08a95
          35478 => x"80", -- $08a96
          35479 => x"80", -- $08a97
          35480 => x"80", -- $08a98
          35481 => x"80", -- $08a99
          35482 => x"80", -- $08a9a
          35483 => x"80", -- $08a9b
          35484 => x"80", -- $08a9c
          35485 => x"80", -- $08a9d
          35486 => x"80", -- $08a9e
          35487 => x"80", -- $08a9f
          35488 => x"80", -- $08aa0
          35489 => x"80", -- $08aa1
          35490 => x"80", -- $08aa2
          35491 => x"80", -- $08aa3
          35492 => x"80", -- $08aa4
          35493 => x"80", -- $08aa5
          35494 => x"80", -- $08aa6
          35495 => x"80", -- $08aa7
          35496 => x"80", -- $08aa8
          35497 => x"80", -- $08aa9
          35498 => x"80", -- $08aaa
          35499 => x"80", -- $08aab
          35500 => x"80", -- $08aac
          35501 => x"80", -- $08aad
          35502 => x"80", -- $08aae
          35503 => x"80", -- $08aaf
          35504 => x"80", -- $08ab0
          35505 => x"80", -- $08ab1
          35506 => x"80", -- $08ab2
          35507 => x"80", -- $08ab3
          35508 => x"80", -- $08ab4
          35509 => x"80", -- $08ab5
          35510 => x"80", -- $08ab6
          35511 => x"80", -- $08ab7
          35512 => x"80", -- $08ab8
          35513 => x"80", -- $08ab9
          35514 => x"80", -- $08aba
          35515 => x"80", -- $08abb
          35516 => x"80", -- $08abc
          35517 => x"80", -- $08abd
          35518 => x"80", -- $08abe
          35519 => x"80", -- $08abf
          35520 => x"80", -- $08ac0
          35521 => x"80", -- $08ac1
          35522 => x"80", -- $08ac2
          35523 => x"80", -- $08ac3
          35524 => x"80", -- $08ac4
          35525 => x"80", -- $08ac5
          35526 => x"80", -- $08ac6
          35527 => x"80", -- $08ac7
          35528 => x"80", -- $08ac8
          35529 => x"80", -- $08ac9
          35530 => x"80", -- $08aca
          35531 => x"80", -- $08acb
          35532 => x"80", -- $08acc
          35533 => x"80", -- $08acd
          35534 => x"80", -- $08ace
          35535 => x"80", -- $08acf
          35536 => x"80", -- $08ad0
          35537 => x"80", -- $08ad1
          35538 => x"80", -- $08ad2
          35539 => x"80", -- $08ad3
          35540 => x"80", -- $08ad4
          35541 => x"80", -- $08ad5
          35542 => x"80", -- $08ad6
          35543 => x"80", -- $08ad7
          35544 => x"80", -- $08ad8
          35545 => x"80", -- $08ad9
          35546 => x"80", -- $08ada
          35547 => x"80", -- $08adb
          35548 => x"80", -- $08adc
          35549 => x"80", -- $08add
          35550 => x"80", -- $08ade
          35551 => x"7f", -- $08adf
          35552 => x"7f", -- $08ae0
          35553 => x"80", -- $08ae1
          35554 => x"80", -- $08ae2
          35555 => x"80", -- $08ae3
          35556 => x"80", -- $08ae4
          35557 => x"80", -- $08ae5
          35558 => x"80", -- $08ae6
          35559 => x"80", -- $08ae7
          35560 => x"80", -- $08ae8
          35561 => x"80", -- $08ae9
          35562 => x"80", -- $08aea
          35563 => x"80", -- $08aeb
          35564 => x"80", -- $08aec
          35565 => x"80", -- $08aed
          35566 => x"80", -- $08aee
          35567 => x"80", -- $08aef
          35568 => x"80", -- $08af0
          35569 => x"80", -- $08af1
          35570 => x"80", -- $08af2
          35571 => x"80", -- $08af3
          35572 => x"80", -- $08af4
          35573 => x"80", -- $08af5
          35574 => x"80", -- $08af6
          35575 => x"80", -- $08af7
          35576 => x"80", -- $08af8
          35577 => x"80", -- $08af9
          35578 => x"80", -- $08afa
          35579 => x"80", -- $08afb
          35580 => x"80", -- $08afc
          35581 => x"80", -- $08afd
          35582 => x"80", -- $08afe
          35583 => x"80", -- $08aff
          35584 => x"80", -- $08b00
          35585 => x"80", -- $08b01
          35586 => x"80", -- $08b02
          35587 => x"80", -- $08b03
          35588 => x"80", -- $08b04
          35589 => x"80", -- $08b05
          35590 => x"80", -- $08b06
          35591 => x"80", -- $08b07
          35592 => x"80", -- $08b08
          35593 => x"80", -- $08b09
          35594 => x"80", -- $08b0a
          35595 => x"80", -- $08b0b
          35596 => x"80", -- $08b0c
          35597 => x"80", -- $08b0d
          35598 => x"80", -- $08b0e
          35599 => x"80", -- $08b0f
          35600 => x"80", -- $08b10
          35601 => x"80", -- $08b11
          35602 => x"80", -- $08b12
          35603 => x"80", -- $08b13
          35604 => x"80", -- $08b14
          35605 => x"80", -- $08b15
          35606 => x"80", -- $08b16
          35607 => x"80", -- $08b17
          35608 => x"80", -- $08b18
          35609 => x"80", -- $08b19
          35610 => x"80", -- $08b1a
          35611 => x"80", -- $08b1b
          35612 => x"80", -- $08b1c
          35613 => x"80", -- $08b1d
          35614 => x"80", -- $08b1e
          35615 => x"80", -- $08b1f
          35616 => x"80", -- $08b20
          35617 => x"80", -- $08b21
          35618 => x"80", -- $08b22
          35619 => x"80", -- $08b23
          35620 => x"80", -- $08b24
          35621 => x"80", -- $08b25
          35622 => x"80", -- $08b26
          35623 => x"80", -- $08b27
          35624 => x"80", -- $08b28
          35625 => x"80", -- $08b29
          35626 => x"80", -- $08b2a
          35627 => x"80", -- $08b2b
          35628 => x"80", -- $08b2c
          35629 => x"80", -- $08b2d
          35630 => x"80", -- $08b2e
          35631 => x"80", -- $08b2f
          35632 => x"80", -- $08b30
          35633 => x"80", -- $08b31
          35634 => x"80", -- $08b32
          35635 => x"80", -- $08b33
          35636 => x"80", -- $08b34
          35637 => x"80", -- $08b35
          35638 => x"80", -- $08b36
          35639 => x"80", -- $08b37
          35640 => x"80", -- $08b38
          35641 => x"7f", -- $08b39
          35642 => x"7f", -- $08b3a
          35643 => x"7f", -- $08b3b
          35644 => x"7f", -- $08b3c
          35645 => x"7f", -- $08b3d
          35646 => x"7f", -- $08b3e
          35647 => x"7f", -- $08b3f
          35648 => x"80", -- $08b40
          35649 => x"80", -- $08b41
          35650 => x"80", -- $08b42
          35651 => x"80", -- $08b43
          35652 => x"80", -- $08b44
          35653 => x"80", -- $08b45
          35654 => x"7f", -- $08b46
          35655 => x"80", -- $08b47
          35656 => x"80", -- $08b48
          35657 => x"80", -- $08b49
          35658 => x"80", -- $08b4a
          35659 => x"80", -- $08b4b
          35660 => x"80", -- $08b4c
          35661 => x"80", -- $08b4d
          35662 => x"80", -- $08b4e
          35663 => x"80", -- $08b4f
          35664 => x"80", -- $08b50
          35665 => x"7f", -- $08b51
          35666 => x"7f", -- $08b52
          35667 => x"7f", -- $08b53
          35668 => x"7f", -- $08b54
          35669 => x"7f", -- $08b55
          35670 => x"7f", -- $08b56
          35671 => x"7f", -- $08b57
          35672 => x"7f", -- $08b58
          35673 => x"7f", -- $08b59
          35674 => x"7f", -- $08b5a
          35675 => x"7f", -- $08b5b
          35676 => x"80", -- $08b5c
          35677 => x"80", -- $08b5d
          35678 => x"80", -- $08b5e
          35679 => x"80", -- $08b5f
          35680 => x"80", -- $08b60
          35681 => x"80", -- $08b61
          35682 => x"80", -- $08b62
          35683 => x"80", -- $08b63
          35684 => x"80", -- $08b64
          35685 => x"7f", -- $08b65
          35686 => x"7f", -- $08b66
          35687 => x"7f", -- $08b67
          35688 => x"80", -- $08b68
          35689 => x"80", -- $08b69
          35690 => x"7f", -- $08b6a
          35691 => x"80", -- $08b6b
          35692 => x"80", -- $08b6c
          35693 => x"7f", -- $08b6d
          35694 => x"7f", -- $08b6e
          35695 => x"7f", -- $08b6f
          35696 => x"7f", -- $08b70
          35697 => x"7f", -- $08b71
          35698 => x"7f", -- $08b72
          35699 => x"7f", -- $08b73
          35700 => x"7f", -- $08b74
          35701 => x"7f", -- $08b75
          35702 => x"7f", -- $08b76
          35703 => x"7f", -- $08b77
          35704 => x"7f", -- $08b78
          35705 => x"7f", -- $08b79
          35706 => x"7f", -- $08b7a
          35707 => x"7f", -- $08b7b
          35708 => x"7f", -- $08b7c
          35709 => x"80", -- $08b7d
          35710 => x"80", -- $08b7e
          35711 => x"80", -- $08b7f
          35712 => x"80", -- $08b80
          35713 => x"80", -- $08b81
          35714 => x"80", -- $08b82
          35715 => x"80", -- $08b83
          35716 => x"80", -- $08b84
          35717 => x"80", -- $08b85
          35718 => x"80", -- $08b86
          35719 => x"80", -- $08b87
          35720 => x"80", -- $08b88
          35721 => x"7f", -- $08b89
          35722 => x"7f", -- $08b8a
          35723 => x"7f", -- $08b8b
          35724 => x"7f", -- $08b8c
          35725 => x"7f", -- $08b8d
          35726 => x"7f", -- $08b8e
          35727 => x"7f", -- $08b8f
          35728 => x"7f", -- $08b90
          35729 => x"7f", -- $08b91
          35730 => x"7f", -- $08b92
          35731 => x"7f", -- $08b93
          35732 => x"7f", -- $08b94
          35733 => x"7f", -- $08b95
          35734 => x"7f", -- $08b96
          35735 => x"7f", -- $08b97
          35736 => x"7f", -- $08b98
          35737 => x"7f", -- $08b99
          35738 => x"7f", -- $08b9a
          35739 => x"7f", -- $08b9b
          35740 => x"7f", -- $08b9c
          35741 => x"80", -- $08b9d
          35742 => x"80", -- $08b9e
          35743 => x"80", -- $08b9f
          35744 => x"80", -- $08ba0
          35745 => x"80", -- $08ba1
          35746 => x"80", -- $08ba2
          35747 => x"80", -- $08ba3
          35748 => x"7f", -- $08ba4
          35749 => x"7f", -- $08ba5
          35750 => x"7f", -- $08ba6
          35751 => x"7f", -- $08ba7
          35752 => x"7f", -- $08ba8
          35753 => x"7f", -- $08ba9
          35754 => x"7f", -- $08baa
          35755 => x"7f", -- $08bab
          35756 => x"7f", -- $08bac
          35757 => x"7f", -- $08bad
          35758 => x"7f", -- $08bae
          35759 => x"7f", -- $08baf
          35760 => x"7f", -- $08bb0
          35761 => x"7f", -- $08bb1
          35762 => x"7f", -- $08bb2
          35763 => x"7f", -- $08bb3
          35764 => x"7f", -- $08bb4
          35765 => x"7f", -- $08bb5
          35766 => x"7f", -- $08bb6
          35767 => x"7f", -- $08bb7
          35768 => x"7f", -- $08bb8
          35769 => x"7f", -- $08bb9
          35770 => x"7f", -- $08bba
          35771 => x"80", -- $08bbb
          35772 => x"7f", -- $08bbc
          35773 => x"7f", -- $08bbd
          35774 => x"7f", -- $08bbe
          35775 => x"80", -- $08bbf
          35776 => x"80", -- $08bc0
          35777 => x"80", -- $08bc1
          35778 => x"80", -- $08bc2
          35779 => x"80", -- $08bc3
          35780 => x"80", -- $08bc4
          35781 => x"80", -- $08bc5
          35782 => x"80", -- $08bc6
          35783 => x"7f", -- $08bc7
          35784 => x"7f", -- $08bc8
          35785 => x"7f", -- $08bc9
          35786 => x"7f", -- $08bca
          35787 => x"7f", -- $08bcb
          35788 => x"7f", -- $08bcc
          35789 => x"7f", -- $08bcd
          35790 => x"7f", -- $08bce
          35791 => x"7f", -- $08bcf
          35792 => x"7f", -- $08bd0
          35793 => x"7f", -- $08bd1
          35794 => x"7f", -- $08bd2
          35795 => x"7f", -- $08bd3
          35796 => x"7f", -- $08bd4
          35797 => x"7f", -- $08bd5
          35798 => x"7f", -- $08bd6
          35799 => x"7f", -- $08bd7
          35800 => x"7f", -- $08bd8
          35801 => x"7f", -- $08bd9
          35802 => x"80", -- $08bda
          35803 => x"80", -- $08bdb
          35804 => x"80", -- $08bdc
          35805 => x"80", -- $08bdd
          35806 => x"80", -- $08bde
          35807 => x"80", -- $08bdf
          35808 => x"80", -- $08be0
          35809 => x"80", -- $08be1
          35810 => x"80", -- $08be2
          35811 => x"80", -- $08be3
          35812 => x"80", -- $08be4
          35813 => x"80", -- $08be5
          35814 => x"7f", -- $08be6
          35815 => x"7f", -- $08be7
          35816 => x"7f", -- $08be8
          35817 => x"7f", -- $08be9
          35818 => x"7f", -- $08bea
          35819 => x"7f", -- $08beb
          35820 => x"7f", -- $08bec
          35821 => x"7f", -- $08bed
          35822 => x"7f", -- $08bee
          35823 => x"7f", -- $08bef
          35824 => x"7f", -- $08bf0
          35825 => x"7f", -- $08bf1
          35826 => x"7f", -- $08bf2
          35827 => x"7f", -- $08bf3
          35828 => x"80", -- $08bf4
          35829 => x"80", -- $08bf5
          35830 => x"80", -- $08bf6
          35831 => x"80", -- $08bf7
          35832 => x"80", -- $08bf8
          35833 => x"80", -- $08bf9
          35834 => x"80", -- $08bfa
          35835 => x"80", -- $08bfb
          35836 => x"80", -- $08bfc
          35837 => x"80", -- $08bfd
          35838 => x"80", -- $08bfe
          35839 => x"80", -- $08bff
          35840 => x"80", -- $08c00
          35841 => x"80", -- $08c01
          35842 => x"80", -- $08c02
          35843 => x"80", -- $08c03
          35844 => x"80", -- $08c04
          35845 => x"80", -- $08c05
          35846 => x"80", -- $08c06
          35847 => x"80", -- $08c07
          35848 => x"80", -- $08c08
          35849 => x"80", -- $08c09
          35850 => x"80", -- $08c0a
          35851 => x"80", -- $08c0b
          35852 => x"80", -- $08c0c
          35853 => x"80", -- $08c0d
          35854 => x"80", -- $08c0e
          35855 => x"80", -- $08c0f
          35856 => x"80", -- $08c10
          35857 => x"80", -- $08c11
          35858 => x"80", -- $08c12
          35859 => x"80", -- $08c13
          35860 => x"80", -- $08c14
          35861 => x"80", -- $08c15
          35862 => x"80", -- $08c16
          35863 => x"80", -- $08c17
          35864 => x"80", -- $08c18
          35865 => x"80", -- $08c19
          35866 => x"80", -- $08c1a
          35867 => x"80", -- $08c1b
          35868 => x"80", -- $08c1c
          35869 => x"80", -- $08c1d
          35870 => x"80", -- $08c1e
          35871 => x"80", -- $08c1f
          35872 => x"80", -- $08c20
          35873 => x"80", -- $08c21
          35874 => x"80", -- $08c22
          35875 => x"80", -- $08c23
          35876 => x"80", -- $08c24
          35877 => x"80", -- $08c25
          35878 => x"80", -- $08c26
          35879 => x"80", -- $08c27
          35880 => x"80", -- $08c28
          35881 => x"80", -- $08c29
          35882 => x"80", -- $08c2a
          35883 => x"80", -- $08c2b
          35884 => x"80", -- $08c2c
          35885 => x"80", -- $08c2d
          35886 => x"80", -- $08c2e
          35887 => x"80", -- $08c2f
          35888 => x"80", -- $08c30
          35889 => x"80", -- $08c31
          35890 => x"80", -- $08c32
          35891 => x"80", -- $08c33
          35892 => x"80", -- $08c34
          35893 => x"80", -- $08c35
          35894 => x"80", -- $08c36
          35895 => x"80", -- $08c37
          35896 => x"80", -- $08c38
          35897 => x"80", -- $08c39
          35898 => x"80", -- $08c3a
          35899 => x"80", -- $08c3b
          35900 => x"80", -- $08c3c
          35901 => x"80", -- $08c3d
          35902 => x"80", -- $08c3e
          35903 => x"80", -- $08c3f
          35904 => x"80", -- $08c40
          35905 => x"80", -- $08c41
          35906 => x"80", -- $08c42
          35907 => x"80", -- $08c43
          35908 => x"80", -- $08c44
          35909 => x"80", -- $08c45
          35910 => x"80", -- $08c46
          35911 => x"80", -- $08c47
          35912 => x"80", -- $08c48
          35913 => x"80", -- $08c49
          35914 => x"80", -- $08c4a
          35915 => x"80", -- $08c4b
          35916 => x"80", -- $08c4c
          35917 => x"80", -- $08c4d
          35918 => x"80", -- $08c4e
          35919 => x"80", -- $08c4f
          35920 => x"80", -- $08c50
          35921 => x"80", -- $08c51
          35922 => x"80", -- $08c52
          35923 => x"80", -- $08c53
          35924 => x"80", -- $08c54
          35925 => x"80", -- $08c55
          35926 => x"80", -- $08c56
          35927 => x"80", -- $08c57
          35928 => x"80", -- $08c58
          35929 => x"80", -- $08c59
          35930 => x"80", -- $08c5a
          35931 => x"80", -- $08c5b
          35932 => x"80", -- $08c5c
          35933 => x"80", -- $08c5d
          35934 => x"80", -- $08c5e
          35935 => x"80", -- $08c5f
          35936 => x"80", -- $08c60
          35937 => x"80", -- $08c61
          35938 => x"80", -- $08c62
          35939 => x"80", -- $08c63
          35940 => x"80", -- $08c64
          35941 => x"80", -- $08c65
          35942 => x"80", -- $08c66
          35943 => x"80", -- $08c67
          35944 => x"80", -- $08c68
          35945 => x"80", -- $08c69
          35946 => x"80", -- $08c6a
          35947 => x"80", -- $08c6b
          35948 => x"80", -- $08c6c
          35949 => x"80", -- $08c6d
          35950 => x"80", -- $08c6e
          35951 => x"80", -- $08c6f
          35952 => x"80", -- $08c70
          35953 => x"80", -- $08c71
          35954 => x"80", -- $08c72
          35955 => x"80", -- $08c73
          35956 => x"80", -- $08c74
          35957 => x"80", -- $08c75
          35958 => x"80", -- $08c76
          35959 => x"80", -- $08c77
          35960 => x"80", -- $08c78
          35961 => x"80", -- $08c79
          35962 => x"80", -- $08c7a
          35963 => x"80", -- $08c7b
          35964 => x"80", -- $08c7c
          35965 => x"80", -- $08c7d
          35966 => x"80", -- $08c7e
          35967 => x"80", -- $08c7f
          35968 => x"80", -- $08c80
          35969 => x"80", -- $08c81
          35970 => x"80", -- $08c82
          35971 => x"80", -- $08c83
          35972 => x"80", -- $08c84
          35973 => x"80", -- $08c85
          35974 => x"80", -- $08c86
          35975 => x"80", -- $08c87
          35976 => x"80", -- $08c88
          35977 => x"80", -- $08c89
          35978 => x"80", -- $08c8a
          35979 => x"80", -- $08c8b
          35980 => x"80", -- $08c8c
          35981 => x"80", -- $08c8d
          35982 => x"80", -- $08c8e
          35983 => x"80", -- $08c8f
          35984 => x"80", -- $08c90
          35985 => x"80", -- $08c91
          35986 => x"80", -- $08c92
          35987 => x"80", -- $08c93
          35988 => x"81", -- $08c94
          35989 => x"81", -- $08c95
          35990 => x"81", -- $08c96
          35991 => x"81", -- $08c97
          35992 => x"81", -- $08c98
          35993 => x"80", -- $08c99
          35994 => x"80", -- $08c9a
          35995 => x"80", -- $08c9b
          35996 => x"80", -- $08c9c
          35997 => x"80", -- $08c9d
          35998 => x"80", -- $08c9e
          35999 => x"80", -- $08c9f
          36000 => x"80", -- $08ca0
          36001 => x"80", -- $08ca1
          36002 => x"80", -- $08ca2
          36003 => x"80", -- $08ca3
          36004 => x"80", -- $08ca4
          36005 => x"80", -- $08ca5
          36006 => x"80", -- $08ca6
          36007 => x"80", -- $08ca7
          36008 => x"80", -- $08ca8
          36009 => x"80", -- $08ca9
          36010 => x"80", -- $08caa
          36011 => x"80", -- $08cab
          36012 => x"80", -- $08cac
          36013 => x"80", -- $08cad
          36014 => x"80", -- $08cae
          36015 => x"81", -- $08caf
          36016 => x"81", -- $08cb0
          36017 => x"81", -- $08cb1
          36018 => x"81", -- $08cb2
          36019 => x"81", -- $08cb3
          36020 => x"81", -- $08cb4
          36021 => x"81", -- $08cb5
          36022 => x"81", -- $08cb6
          36023 => x"81", -- $08cb7
          36024 => x"81", -- $08cb8
          36025 => x"81", -- $08cb9
          36026 => x"81", -- $08cba
          36027 => x"81", -- $08cbb
          36028 => x"81", -- $08cbc
          36029 => x"81", -- $08cbd
          36030 => x"81", -- $08cbe
          36031 => x"81", -- $08cbf
          36032 => x"80", -- $08cc0
          36033 => x"80", -- $08cc1
          36034 => x"80", -- $08cc2
          36035 => x"80", -- $08cc3
          36036 => x"80", -- $08cc4
          36037 => x"80", -- $08cc5
          36038 => x"80", -- $08cc6
          36039 => x"80", -- $08cc7
          36040 => x"80", -- $08cc8
          36041 => x"80", -- $08cc9
          36042 => x"81", -- $08cca
          36043 => x"81", -- $08ccb
          36044 => x"81", -- $08ccc
          36045 => x"81", -- $08ccd
          36046 => x"81", -- $08cce
          36047 => x"81", -- $08ccf
          36048 => x"81", -- $08cd0
          36049 => x"81", -- $08cd1
          36050 => x"81", -- $08cd2
          36051 => x"81", -- $08cd3
          36052 => x"81", -- $08cd4
          36053 => x"81", -- $08cd5
          36054 => x"81", -- $08cd6
          36055 => x"81", -- $08cd7
          36056 => x"81", -- $08cd8
          36057 => x"81", -- $08cd9
          36058 => x"81", -- $08cda
          36059 => x"81", -- $08cdb
          36060 => x"81", -- $08cdc
          36061 => x"81", -- $08cdd
          36062 => x"81", -- $08cde
          36063 => x"81", -- $08cdf
          36064 => x"80", -- $08ce0
          36065 => x"80", -- $08ce1
          36066 => x"80", -- $08ce2
          36067 => x"80", -- $08ce3
          36068 => x"80", -- $08ce4
          36069 => x"80", -- $08ce5
          36070 => x"80", -- $08ce6
          36071 => x"80", -- $08ce7
          36072 => x"80", -- $08ce8
          36073 => x"80", -- $08ce9
          36074 => x"80", -- $08cea
          36075 => x"81", -- $08ceb
          36076 => x"81", -- $08cec
          36077 => x"81", -- $08ced
          36078 => x"81", -- $08cee
          36079 => x"81", -- $08cef
          36080 => x"81", -- $08cf0
          36081 => x"81", -- $08cf1
          36082 => x"81", -- $08cf2
          36083 => x"81", -- $08cf3
          36084 => x"81", -- $08cf4
          36085 => x"81", -- $08cf5
          36086 => x"81", -- $08cf6
          36087 => x"81", -- $08cf7
          36088 => x"81", -- $08cf8
          36089 => x"81", -- $08cf9
          36090 => x"81", -- $08cfa
          36091 => x"81", -- $08cfb
          36092 => x"81", -- $08cfc
          36093 => x"81", -- $08cfd
          36094 => x"81", -- $08cfe
          36095 => x"80", -- $08cff
          36096 => x"80", -- $08d00
          36097 => x"80", -- $08d01
          36098 => x"80", -- $08d02
          36099 => x"80", -- $08d03
          36100 => x"80", -- $08d04
          36101 => x"80", -- $08d05
          36102 => x"80", -- $08d06
          36103 => x"80", -- $08d07
          36104 => x"80", -- $08d08
          36105 => x"80", -- $08d09
          36106 => x"80", -- $08d0a
          36107 => x"81", -- $08d0b
          36108 => x"81", -- $08d0c
          36109 => x"81", -- $08d0d
          36110 => x"81", -- $08d0e
          36111 => x"81", -- $08d0f
          36112 => x"81", -- $08d10
          36113 => x"81", -- $08d11
          36114 => x"81", -- $08d12
          36115 => x"81", -- $08d13
          36116 => x"81", -- $08d14
          36117 => x"81", -- $08d15
          36118 => x"81", -- $08d16
          36119 => x"81", -- $08d17
          36120 => x"81", -- $08d18
          36121 => x"81", -- $08d19
          36122 => x"80", -- $08d1a
          36123 => x"80", -- $08d1b
          36124 => x"80", -- $08d1c
          36125 => x"80", -- $08d1d
          36126 => x"80", -- $08d1e
          36127 => x"80", -- $08d1f
          36128 => x"80", -- $08d20
          36129 => x"80", -- $08d21
          36130 => x"80", -- $08d22
          36131 => x"80", -- $08d23
          36132 => x"80", -- $08d24
          36133 => x"80", -- $08d25
          36134 => x"80", -- $08d26
          36135 => x"80", -- $08d27
          36136 => x"80", -- $08d28
          36137 => x"80", -- $08d29
          36138 => x"80", -- $08d2a
          36139 => x"80", -- $08d2b
          36140 => x"80", -- $08d2c
          36141 => x"80", -- $08d2d
          36142 => x"80", -- $08d2e
          36143 => x"80", -- $08d2f
          36144 => x"80", -- $08d30
          36145 => x"80", -- $08d31
          36146 => x"80", -- $08d32
          36147 => x"80", -- $08d33
          36148 => x"80", -- $08d34
          36149 => x"80", -- $08d35
          36150 => x"80", -- $08d36
          36151 => x"80", -- $08d37
          36152 => x"80", -- $08d38
          36153 => x"80", -- $08d39
          36154 => x"80", -- $08d3a
          36155 => x"80", -- $08d3b
          36156 => x"80", -- $08d3c
          36157 => x"80", -- $08d3d
          36158 => x"80", -- $08d3e
          36159 => x"80", -- $08d3f
          36160 => x"80", -- $08d40
          36161 => x"80", -- $08d41
          36162 => x"80", -- $08d42
          36163 => x"80", -- $08d43
          36164 => x"80", -- $08d44
          36165 => x"80", -- $08d45
          36166 => x"80", -- $08d46
          36167 => x"80", -- $08d47
          36168 => x"80", -- $08d48
          36169 => x"80", -- $08d49
          36170 => x"80", -- $08d4a
          36171 => x"80", -- $08d4b
          36172 => x"80", -- $08d4c
          36173 => x"80", -- $08d4d
          36174 => x"80", -- $08d4e
          36175 => x"80", -- $08d4f
          36176 => x"80", -- $08d50
          36177 => x"80", -- $08d51
          36178 => x"80", -- $08d52
          36179 => x"80", -- $08d53
          36180 => x"80", -- $08d54
          36181 => x"80", -- $08d55
          36182 => x"80", -- $08d56
          36183 => x"80", -- $08d57
          36184 => x"80", -- $08d58
          36185 => x"80", -- $08d59
          36186 => x"80", -- $08d5a
          36187 => x"80", -- $08d5b
          36188 => x"80", -- $08d5c
          36189 => x"80", -- $08d5d
          36190 => x"80", -- $08d5e
          36191 => x"80", -- $08d5f
          36192 => x"80", -- $08d60
          36193 => x"80", -- $08d61
          36194 => x"80", -- $08d62
          36195 => x"80", -- $08d63
          36196 => x"80", -- $08d64
          36197 => x"80", -- $08d65
          36198 => x"80", -- $08d66
          36199 => x"80", -- $08d67
          36200 => x"80", -- $08d68
          36201 => x"80", -- $08d69
          36202 => x"80", -- $08d6a
          36203 => x"80", -- $08d6b
          36204 => x"80", -- $08d6c
          36205 => x"80", -- $08d6d
          36206 => x"80", -- $08d6e
          36207 => x"80", -- $08d6f
          36208 => x"81", -- $08d70
          36209 => x"81", -- $08d71
          36210 => x"81", -- $08d72
          36211 => x"81", -- $08d73
          36212 => x"80", -- $08d74
          36213 => x"80", -- $08d75
          36214 => x"80", -- $08d76
          36215 => x"80", -- $08d77
          36216 => x"80", -- $08d78
          36217 => x"80", -- $08d79
          36218 => x"80", -- $08d7a
          36219 => x"80", -- $08d7b
          36220 => x"80", -- $08d7c
          36221 => x"80", -- $08d7d
          36222 => x"80", -- $08d7e
          36223 => x"80", -- $08d7f
          36224 => x"80", -- $08d80
          36225 => x"80", -- $08d81
          36226 => x"80", -- $08d82
          36227 => x"80", -- $08d83
          36228 => x"80", -- $08d84
          36229 => x"80", -- $08d85
          36230 => x"80", -- $08d86
          36231 => x"80", -- $08d87
          36232 => x"80", -- $08d88
          36233 => x"80", -- $08d89
          36234 => x"80", -- $08d8a
          36235 => x"80", -- $08d8b
          36236 => x"81", -- $08d8c
          36237 => x"81", -- $08d8d
          36238 => x"81", -- $08d8e
          36239 => x"81", -- $08d8f
          36240 => x"81", -- $08d90
          36241 => x"81", -- $08d91
          36242 => x"80", -- $08d92
          36243 => x"80", -- $08d93
          36244 => x"80", -- $08d94
          36245 => x"80", -- $08d95
          36246 => x"80", -- $08d96
          36247 => x"80", -- $08d97
          36248 => x"80", -- $08d98
          36249 => x"80", -- $08d99
          36250 => x"80", -- $08d9a
          36251 => x"80", -- $08d9b
          36252 => x"80", -- $08d9c
          36253 => x"80", -- $08d9d
          36254 => x"80", -- $08d9e
          36255 => x"80", -- $08d9f
          36256 => x"80", -- $08da0
          36257 => x"80", -- $08da1
          36258 => x"80", -- $08da2
          36259 => x"80", -- $08da3
          36260 => x"80", -- $08da4
          36261 => x"80", -- $08da5
          36262 => x"80", -- $08da6
          36263 => x"80", -- $08da7
          36264 => x"80", -- $08da8
          36265 => x"80", -- $08da9
          36266 => x"80", -- $08daa
          36267 => x"80", -- $08dab
          36268 => x"80", -- $08dac
          36269 => x"80", -- $08dad
          36270 => x"81", -- $08dae
          36271 => x"80", -- $08daf
          36272 => x"80", -- $08db0
          36273 => x"80", -- $08db1
          36274 => x"80", -- $08db2
          36275 => x"80", -- $08db3
          36276 => x"80", -- $08db4
          36277 => x"80", -- $08db5
          36278 => x"80", -- $08db6
          36279 => x"80", -- $08db7
          36280 => x"80", -- $08db8
          36281 => x"80", -- $08db9
          36282 => x"80", -- $08dba
          36283 => x"80", -- $08dbb
          36284 => x"80", -- $08dbc
          36285 => x"80", -- $08dbd
          36286 => x"80", -- $08dbe
          36287 => x"80", -- $08dbf
          36288 => x"80", -- $08dc0
          36289 => x"80", -- $08dc1
          36290 => x"80", -- $08dc2
          36291 => x"80", -- $08dc3
          36292 => x"80", -- $08dc4
          36293 => x"80", -- $08dc5
          36294 => x"80", -- $08dc6
          36295 => x"80", -- $08dc7
          36296 => x"80", -- $08dc8
          36297 => x"80", -- $08dc9
          36298 => x"80", -- $08dca
          36299 => x"80", -- $08dcb
          36300 => x"80", -- $08dcc
          36301 => x"80", -- $08dcd
          36302 => x"80", -- $08dce
          36303 => x"80", -- $08dcf
          36304 => x"80", -- $08dd0
          36305 => x"80", -- $08dd1
          36306 => x"80", -- $08dd2
          36307 => x"80", -- $08dd3
          36308 => x"80", -- $08dd4
          36309 => x"80", -- $08dd5
          36310 => x"80", -- $08dd6
          36311 => x"80", -- $08dd7
          36312 => x"80", -- $08dd8
          36313 => x"80", -- $08dd9
          36314 => x"80", -- $08dda
          36315 => x"7f", -- $08ddb
          36316 => x"7f", -- $08ddc
          36317 => x"7f", -- $08ddd
          36318 => x"7f", -- $08dde
          36319 => x"7f", -- $08ddf
          36320 => x"80", -- $08de0
          36321 => x"80", -- $08de1
          36322 => x"80", -- $08de2
          36323 => x"80", -- $08de3
          36324 => x"80", -- $08de4
          36325 => x"80", -- $08de5
          36326 => x"80", -- $08de6
          36327 => x"80", -- $08de7
          36328 => x"80", -- $08de8
          36329 => x"80", -- $08de9
          36330 => x"80", -- $08dea
          36331 => x"80", -- $08deb
          36332 => x"80", -- $08dec
          36333 => x"80", -- $08ded
          36334 => x"80", -- $08dee
          36335 => x"80", -- $08def
          36336 => x"80", -- $08df0
          36337 => x"80", -- $08df1
          36338 => x"80", -- $08df2
          36339 => x"80", -- $08df3
          36340 => x"80", -- $08df4
          36341 => x"80", -- $08df5
          36342 => x"80", -- $08df6
          36343 => x"7f", -- $08df7
          36344 => x"7f", -- $08df8
          36345 => x"7f", -- $08df9
          36346 => x"7f", -- $08dfa
          36347 => x"7f", -- $08dfb
          36348 => x"7f", -- $08dfc
          36349 => x"7f", -- $08dfd
          36350 => x"7f", -- $08dfe
          36351 => x"7f", -- $08dff
          36352 => x"7f", -- $08e00
          36353 => x"7f", -- $08e01
          36354 => x"80", -- $08e02
          36355 => x"80", -- $08e03
          36356 => x"80", -- $08e04
          36357 => x"80", -- $08e05
          36358 => x"80", -- $08e06
          36359 => x"80", -- $08e07
          36360 => x"80", -- $08e08
          36361 => x"80", -- $08e09
          36362 => x"80", -- $08e0a
          36363 => x"80", -- $08e0b
          36364 => x"80", -- $08e0c
          36365 => x"80", -- $08e0d
          36366 => x"80", -- $08e0e
          36367 => x"80", -- $08e0f
          36368 => x"80", -- $08e10
          36369 => x"80", -- $08e11
          36370 => x"80", -- $08e12
          36371 => x"80", -- $08e13
          36372 => x"7f", -- $08e14
          36373 => x"7f", -- $08e15
          36374 => x"7f", -- $08e16
          36375 => x"7f", -- $08e17
          36376 => x"7f", -- $08e18
          36377 => x"7e", -- $08e19
          36378 => x"7e", -- $08e1a
          36379 => x"7e", -- $08e1b
          36380 => x"7e", -- $08e1c
          36381 => x"7f", -- $08e1d
          36382 => x"7f", -- $08e1e
          36383 => x"7f", -- $08e1f
          36384 => x"7f", -- $08e20
          36385 => x"7f", -- $08e21
          36386 => x"7f", -- $08e22
          36387 => x"80", -- $08e23
          36388 => x"80", -- $08e24
          36389 => x"80", -- $08e25
          36390 => x"80", -- $08e26
          36391 => x"80", -- $08e27
          36392 => x"80", -- $08e28
          36393 => x"80", -- $08e29
          36394 => x"80", -- $08e2a
          36395 => x"80", -- $08e2b
          36396 => x"80", -- $08e2c
          36397 => x"80", -- $08e2d
          36398 => x"80", -- $08e2e
          36399 => x"80", -- $08e2f
          36400 => x"80", -- $08e30
          36401 => x"7f", -- $08e31
          36402 => x"7f", -- $08e32
          36403 => x"7f", -- $08e33
          36404 => x"7f", -- $08e34
          36405 => x"7f", -- $08e35
          36406 => x"7f", -- $08e36
          36407 => x"7e", -- $08e37
          36408 => x"7e", -- $08e38
          36409 => x"7e", -- $08e39
          36410 => x"7e", -- $08e3a
          36411 => x"7e", -- $08e3b
          36412 => x"7e", -- $08e3c
          36413 => x"7e", -- $08e3d
          36414 => x"7f", -- $08e3e
          36415 => x"7f", -- $08e3f
          36416 => x"7f", -- $08e40
          36417 => x"7f", -- $08e41
          36418 => x"7f", -- $08e42
          36419 => x"7f", -- $08e43
          36420 => x"80", -- $08e44
          36421 => x"80", -- $08e45
          36422 => x"80", -- $08e46
          36423 => x"80", -- $08e47
          36424 => x"80", -- $08e48
          36425 => x"80", -- $08e49
          36426 => x"80", -- $08e4a
          36427 => x"80", -- $08e4b
          36428 => x"80", -- $08e4c
          36429 => x"80", -- $08e4d
          36430 => x"80", -- $08e4e
          36431 => x"7f", -- $08e4f
          36432 => x"7f", -- $08e50
          36433 => x"7f", -- $08e51
          36434 => x"7f", -- $08e52
          36435 => x"7f", -- $08e53
          36436 => x"7e", -- $08e54
          36437 => x"7e", -- $08e55
          36438 => x"7e", -- $08e56
          36439 => x"7e", -- $08e57
          36440 => x"7e", -- $08e58
          36441 => x"7e", -- $08e59
          36442 => x"7e", -- $08e5a
          36443 => x"7e", -- $08e5b
          36444 => x"7e", -- $08e5c
          36445 => x"7f", -- $08e5d
          36446 => x"7f", -- $08e5e
          36447 => x"7f", -- $08e5f
          36448 => x"7f", -- $08e60
          36449 => x"7f", -- $08e61
          36450 => x"80", -- $08e62
          36451 => x"80", -- $08e63
          36452 => x"80", -- $08e64
          36453 => x"80", -- $08e65
          36454 => x"80", -- $08e66
          36455 => x"80", -- $08e67
          36456 => x"80", -- $08e68
          36457 => x"80", -- $08e69
          36458 => x"80", -- $08e6a
          36459 => x"80", -- $08e6b
          36460 => x"80", -- $08e6c
          36461 => x"80", -- $08e6d
          36462 => x"80", -- $08e6e
          36463 => x"80", -- $08e6f
          36464 => x"7f", -- $08e70
          36465 => x"7f", -- $08e71
          36466 => x"7f", -- $08e72
          36467 => x"7f", -- $08e73
          36468 => x"7f", -- $08e74
          36469 => x"7f", -- $08e75
          36470 => x"7f", -- $08e76
          36471 => x"7f", -- $08e77
          36472 => x"7f", -- $08e78
          36473 => x"7f", -- $08e79
          36474 => x"7f", -- $08e7a
          36475 => x"7f", -- $08e7b
          36476 => x"7f", -- $08e7c
          36477 => x"7f", -- $08e7d
          36478 => x"80", -- $08e7e
          36479 => x"80", -- $08e7f
          36480 => x"80", -- $08e80
          36481 => x"80", -- $08e81
          36482 => x"80", -- $08e82
          36483 => x"80", -- $08e83
          36484 => x"80", -- $08e84
          36485 => x"80", -- $08e85
          36486 => x"80", -- $08e86
          36487 => x"80", -- $08e87
          36488 => x"80", -- $08e88
          36489 => x"80", -- $08e89
          36490 => x"80", -- $08e8a
          36491 => x"80", -- $08e8b
          36492 => x"80", -- $08e8c
          36493 => x"80", -- $08e8d
          36494 => x"80", -- $08e8e
          36495 => x"80", -- $08e8f
          36496 => x"80", -- $08e90
          36497 => x"80", -- $08e91
          36498 => x"80", -- $08e92
          36499 => x"80", -- $08e93
          36500 => x"80", -- $08e94
          36501 => x"7f", -- $08e95
          36502 => x"7f", -- $08e96
          36503 => x"7f", -- $08e97
          36504 => x"7f", -- $08e98
          36505 => x"7f", -- $08e99
          36506 => x"80", -- $08e9a
          36507 => x"80", -- $08e9b
          36508 => x"80", -- $08e9c
          36509 => x"80", -- $08e9d
          36510 => x"80", -- $08e9e
          36511 => x"80", -- $08e9f
          36512 => x"80", -- $08ea0
          36513 => x"80", -- $08ea1
          36514 => x"80", -- $08ea2
          36515 => x"80", -- $08ea3
          36516 => x"80", -- $08ea4
          36517 => x"80", -- $08ea5
          36518 => x"80", -- $08ea6
          36519 => x"80", -- $08ea7
          36520 => x"80", -- $08ea8
          36521 => x"80", -- $08ea9
          36522 => x"80", -- $08eaa
          36523 => x"80", -- $08eab
          36524 => x"80", -- $08eac
          36525 => x"80", -- $08ead
          36526 => x"80", -- $08eae
          36527 => x"80", -- $08eaf
          36528 => x"80", -- $08eb0
          36529 => x"80", -- $08eb1
          36530 => x"80", -- $08eb2
          36531 => x"80", -- $08eb3
          36532 => x"80", -- $08eb4
          36533 => x"80", -- $08eb5
          36534 => x"80", -- $08eb6
          36535 => x"80", -- $08eb7
          36536 => x"80", -- $08eb8
          36537 => x"80", -- $08eb9
          36538 => x"80", -- $08eba
          36539 => x"80", -- $08ebb
          36540 => x"80", -- $08ebc
          36541 => x"80", -- $08ebd
          36542 => x"80", -- $08ebe
          36543 => x"80", -- $08ebf
          36544 => x"80", -- $08ec0
          36545 => x"80", -- $08ec1
          36546 => x"80", -- $08ec2
          36547 => x"80", -- $08ec3
          36548 => x"80", -- $08ec4
          36549 => x"80", -- $08ec5
          36550 => x"80", -- $08ec6
          36551 => x"80", -- $08ec7
          36552 => x"80", -- $08ec8
          36553 => x"80", -- $08ec9
          36554 => x"80", -- $08eca
          36555 => x"80", -- $08ecb
          36556 => x"80", -- $08ecc
          36557 => x"80", -- $08ecd
          36558 => x"80", -- $08ece
          36559 => x"80", -- $08ecf
          36560 => x"80", -- $08ed0
          36561 => x"80", -- $08ed1
          36562 => x"80", -- $08ed2
          36563 => x"80", -- $08ed3
          36564 => x"80", -- $08ed4
          36565 => x"7f", -- $08ed5
          36566 => x"7f", -- $08ed6
          36567 => x"80", -- $08ed7
          36568 => x"7f", -- $08ed8
          36569 => x"80", -- $08ed9
          36570 => x"80", -- $08eda
          36571 => x"80", -- $08edb
          36572 => x"80", -- $08edc
          36573 => x"80", -- $08edd
          36574 => x"80", -- $08ede
          36575 => x"80", -- $08edf
          36576 => x"80", -- $08ee0
          36577 => x"80", -- $08ee1
          36578 => x"80", -- $08ee2
          36579 => x"80", -- $08ee3
          36580 => x"80", -- $08ee4
          36581 => x"80", -- $08ee5
          36582 => x"80", -- $08ee6
          36583 => x"80", -- $08ee7
          36584 => x"80", -- $08ee8
          36585 => x"80", -- $08ee9
          36586 => x"80", -- $08eea
          36587 => x"80", -- $08eeb
          36588 => x"80", -- $08eec
          36589 => x"80", -- $08eed
          36590 => x"80", -- $08eee
          36591 => x"80", -- $08eef
          36592 => x"7f", -- $08ef0
          36593 => x"7f", -- $08ef1
          36594 => x"7f", -- $08ef2
          36595 => x"7f", -- $08ef3
          36596 => x"7f", -- $08ef4
          36597 => x"7f", -- $08ef5
          36598 => x"7f", -- $08ef6
          36599 => x"7f", -- $08ef7
          36600 => x"7f", -- $08ef8
          36601 => x"80", -- $08ef9
          36602 => x"80", -- $08efa
          36603 => x"80", -- $08efb
          36604 => x"80", -- $08efc
          36605 => x"80", -- $08efd
          36606 => x"80", -- $08efe
          36607 => x"80", -- $08eff
          36608 => x"80", -- $08f00
          36609 => x"80", -- $08f01
          36610 => x"80", -- $08f02
          36611 => x"80", -- $08f03
          36612 => x"80", -- $08f04
          36613 => x"80", -- $08f05
          36614 => x"80", -- $08f06
          36615 => x"80", -- $08f07
          36616 => x"80", -- $08f08
          36617 => x"80", -- $08f09
          36618 => x"80", -- $08f0a
          36619 => x"80", -- $08f0b
          36620 => x"80", -- $08f0c
          36621 => x"80", -- $08f0d
          36622 => x"7f", -- $08f0e
          36623 => x"7f", -- $08f0f
          36624 => x"7f", -- $08f10
          36625 => x"7f", -- $08f11
          36626 => x"7f", -- $08f12
          36627 => x"7f", -- $08f13
          36628 => x"7f", -- $08f14
          36629 => x"7f", -- $08f15
          36630 => x"7f", -- $08f16
          36631 => x"7f", -- $08f17
          36632 => x"7f", -- $08f18
          36633 => x"80", -- $08f19
          36634 => x"80", -- $08f1a
          36635 => x"80", -- $08f1b
          36636 => x"80", -- $08f1c
          36637 => x"80", -- $08f1d
          36638 => x"80", -- $08f1e
          36639 => x"80", -- $08f1f
          36640 => x"80", -- $08f20
          36641 => x"80", -- $08f21
          36642 => x"80", -- $08f22
          36643 => x"80", -- $08f23
          36644 => x"80", -- $08f24
          36645 => x"80", -- $08f25
          36646 => x"80", -- $08f26
          36647 => x"80", -- $08f27
          36648 => x"80", -- $08f28
          36649 => x"80", -- $08f29
          36650 => x"80", -- $08f2a
          36651 => x"80", -- $08f2b
          36652 => x"80", -- $08f2c
          36653 => x"80", -- $08f2d
          36654 => x"80", -- $08f2e
          36655 => x"80", -- $08f2f
          36656 => x"80", -- $08f30
          36657 => x"80", -- $08f31
          36658 => x"80", -- $08f32
          36659 => x"80", -- $08f33
          36660 => x"80", -- $08f34
          36661 => x"80", -- $08f35
          36662 => x"80", -- $08f36
          36663 => x"80", -- $08f37
          36664 => x"80", -- $08f38
          36665 => x"80", -- $08f39
          36666 => x"80", -- $08f3a
          36667 => x"80", -- $08f3b
          36668 => x"80", -- $08f3c
          36669 => x"80", -- $08f3d
          36670 => x"81", -- $08f3e
          36671 => x"81", -- $08f3f
          36672 => x"81", -- $08f40
          36673 => x"81", -- $08f41
          36674 => x"81", -- $08f42
          36675 => x"81", -- $08f43
          36676 => x"81", -- $08f44
          36677 => x"81", -- $08f45
          36678 => x"81", -- $08f46
          36679 => x"81", -- $08f47
          36680 => x"81", -- $08f48
          36681 => x"81", -- $08f49
          36682 => x"80", -- $08f4a
          36683 => x"80", -- $08f4b
          36684 => x"80", -- $08f4c
          36685 => x"80", -- $08f4d
          36686 => x"80", -- $08f4e
          36687 => x"80", -- $08f4f
          36688 => x"80", -- $08f50
          36689 => x"80", -- $08f51
          36690 => x"80", -- $08f52
          36691 => x"80", -- $08f53
          36692 => x"80", -- $08f54
          36693 => x"80", -- $08f55
          36694 => x"80", -- $08f56
          36695 => x"80", -- $08f57
          36696 => x"80", -- $08f58
          36697 => x"80", -- $08f59
          36698 => x"80", -- $08f5a
          36699 => x"81", -- $08f5b
          36700 => x"81", -- $08f5c
          36701 => x"81", -- $08f5d
          36702 => x"81", -- $08f5e
          36703 => x"81", -- $08f5f
          36704 => x"81", -- $08f60
          36705 => x"81", -- $08f61
          36706 => x"82", -- $08f62
          36707 => x"82", -- $08f63
          36708 => x"82", -- $08f64
          36709 => x"81", -- $08f65
          36710 => x"81", -- $08f66
          36711 => x"81", -- $08f67
          36712 => x"81", -- $08f68
          36713 => x"81", -- $08f69
          36714 => x"81", -- $08f6a
          36715 => x"80", -- $08f6b
          36716 => x"80", -- $08f6c
          36717 => x"80", -- $08f6d
          36718 => x"80", -- $08f6e
          36719 => x"80", -- $08f6f
          36720 => x"80", -- $08f70
          36721 => x"80", -- $08f71
          36722 => x"80", -- $08f72
          36723 => x"80", -- $08f73
          36724 => x"80", -- $08f74
          36725 => x"80", -- $08f75
          36726 => x"80", -- $08f76
          36727 => x"80", -- $08f77
          36728 => x"80", -- $08f78
          36729 => x"80", -- $08f79
          36730 => x"80", -- $08f7a
          36731 => x"81", -- $08f7b
          36732 => x"81", -- $08f7c
          36733 => x"81", -- $08f7d
          36734 => x"81", -- $08f7e
          36735 => x"81", -- $08f7f
          36736 => x"81", -- $08f80
          36737 => x"81", -- $08f81
          36738 => x"81", -- $08f82
          36739 => x"81", -- $08f83
          36740 => x"81", -- $08f84
          36741 => x"81", -- $08f85
          36742 => x"81", -- $08f86
          36743 => x"81", -- $08f87
          36744 => x"81", -- $08f88
          36745 => x"81", -- $08f89
          36746 => x"81", -- $08f8a
          36747 => x"80", -- $08f8b
          36748 => x"80", -- $08f8c
          36749 => x"80", -- $08f8d
          36750 => x"80", -- $08f8e
          36751 => x"80", -- $08f8f
          36752 => x"80", -- $08f90
          36753 => x"80", -- $08f91
          36754 => x"80", -- $08f92
          36755 => x"80", -- $08f93
          36756 => x"80", -- $08f94
          36757 => x"80", -- $08f95
          36758 => x"80", -- $08f96
          36759 => x"80", -- $08f97
          36760 => x"80", -- $08f98
          36761 => x"80", -- $08f99
          36762 => x"80", -- $08f9a
          36763 => x"80", -- $08f9b
          36764 => x"80", -- $08f9c
          36765 => x"80", -- $08f9d
          36766 => x"80", -- $08f9e
          36767 => x"80", -- $08f9f
          36768 => x"80", -- $08fa0
          36769 => x"80", -- $08fa1
          36770 => x"80", -- $08fa2
          36771 => x"81", -- $08fa3
          36772 => x"81", -- $08fa4
          36773 => x"81", -- $08fa5
          36774 => x"80", -- $08fa6
          36775 => x"80", -- $08fa7
          36776 => x"80", -- $08fa8
          36777 => x"80", -- $08fa9
          36778 => x"80", -- $08faa
          36779 => x"80", -- $08fab
          36780 => x"80", -- $08fac
          36781 => x"80", -- $08fad
          36782 => x"80", -- $08fae
          36783 => x"80", -- $08faf
          36784 => x"80", -- $08fb0
          36785 => x"80", -- $08fb1
          36786 => x"80", -- $08fb2
          36787 => x"80", -- $08fb3
          36788 => x"80", -- $08fb4
          36789 => x"80", -- $08fb5
          36790 => x"80", -- $08fb6
          36791 => x"80", -- $08fb7
          36792 => x"80", -- $08fb8
          36793 => x"80", -- $08fb9
          36794 => x"80", -- $08fba
          36795 => x"80", -- $08fbb
          36796 => x"80", -- $08fbc
          36797 => x"80", -- $08fbd
          36798 => x"80", -- $08fbe
          36799 => x"80", -- $08fbf
          36800 => x"80", -- $08fc0
          36801 => x"80", -- $08fc1
          36802 => x"80", -- $08fc2
          36803 => x"80", -- $08fc3
          36804 => x"80", -- $08fc4
          36805 => x"80", -- $08fc5
          36806 => x"80", -- $08fc6
          36807 => x"80", -- $08fc7
          36808 => x"80", -- $08fc8
          36809 => x"80", -- $08fc9
          36810 => x"80", -- $08fca
          36811 => x"80", -- $08fcb
          36812 => x"80", -- $08fcc
          36813 => x"80", -- $08fcd
          36814 => x"80", -- $08fce
          36815 => x"80", -- $08fcf
          36816 => x"80", -- $08fd0
          36817 => x"80", -- $08fd1
          36818 => x"80", -- $08fd2
          36819 => x"80", -- $08fd3
          36820 => x"80", -- $08fd4
          36821 => x"80", -- $08fd5
          36822 => x"80", -- $08fd6
          36823 => x"80", -- $08fd7
          36824 => x"80", -- $08fd8
          36825 => x"80", -- $08fd9
          36826 => x"80", -- $08fda
          36827 => x"80", -- $08fdb
          36828 => x"80", -- $08fdc
          36829 => x"80", -- $08fdd
          36830 => x"80", -- $08fde
          36831 => x"80", -- $08fdf
          36832 => x"80", -- $08fe0
          36833 => x"80", -- $08fe1
          36834 => x"80", -- $08fe2
          36835 => x"80", -- $08fe3
          36836 => x"80", -- $08fe4
          36837 => x"80", -- $08fe5
          36838 => x"80", -- $08fe6
          36839 => x"80", -- $08fe7
          36840 => x"80", -- $08fe8
          36841 => x"80", -- $08fe9
          36842 => x"80", -- $08fea
          36843 => x"80", -- $08feb
          36844 => x"80", -- $08fec
          36845 => x"80", -- $08fed
          36846 => x"80", -- $08fee
          36847 => x"80", -- $08fef
          36848 => x"80", -- $08ff0
          36849 => x"80", -- $08ff1
          36850 => x"80", -- $08ff2
          36851 => x"80", -- $08ff3
          36852 => x"80", -- $08ff4
          36853 => x"80", -- $08ff5
          36854 => x"80", -- $08ff6
          36855 => x"80", -- $08ff7
          36856 => x"80", -- $08ff8
          36857 => x"80", -- $08ff9
          36858 => x"80", -- $08ffa
          36859 => x"80", -- $08ffb
          36860 => x"80", -- $08ffc
          36861 => x"80", -- $08ffd
          36862 => x"80", -- $08ffe
          36863 => x"80", -- $08fff
          36864 => x"80", -- $09000
          36865 => x"80", -- $09001
          36866 => x"80", -- $09002
          36867 => x"80", -- $09003
          36868 => x"80", -- $09004
          36869 => x"80", -- $09005
          36870 => x"80", -- $09006
          36871 => x"80", -- $09007
          36872 => x"80", -- $09008
          36873 => x"80", -- $09009
          36874 => x"80", -- $0900a
          36875 => x"80", -- $0900b
          36876 => x"80", -- $0900c
          36877 => x"80", -- $0900d
          36878 => x"80", -- $0900e
          36879 => x"80", -- $0900f
          36880 => x"80", -- $09010
          36881 => x"80", -- $09011
          36882 => x"80", -- $09012
          36883 => x"80", -- $09013
          36884 => x"80", -- $09014
          36885 => x"80", -- $09015
          36886 => x"80", -- $09016
          36887 => x"80", -- $09017
          36888 => x"80", -- $09018
          36889 => x"80", -- $09019
          36890 => x"80", -- $0901a
          36891 => x"80", -- $0901b
          36892 => x"80", -- $0901c
          36893 => x"80", -- $0901d
          36894 => x"80", -- $0901e
          36895 => x"80", -- $0901f
          36896 => x"80", -- $09020
          36897 => x"80", -- $09021
          36898 => x"80", -- $09022
          36899 => x"80", -- $09023
          36900 => x"80", -- $09024
          36901 => x"80", -- $09025
          36902 => x"80", -- $09026
          36903 => x"80", -- $09027
          36904 => x"80", -- $09028
          36905 => x"80", -- $09029
          36906 => x"80", -- $0902a
          36907 => x"80", -- $0902b
          36908 => x"80", -- $0902c
          36909 => x"80", -- $0902d
          36910 => x"80", -- $0902e
          36911 => x"80", -- $0902f
          36912 => x"80", -- $09030
          36913 => x"80", -- $09031
          36914 => x"80", -- $09032
          36915 => x"80", -- $09033
          36916 => x"80", -- $09034
          36917 => x"80", -- $09035
          36918 => x"80", -- $09036
          36919 => x"80", -- $09037
          36920 => x"80", -- $09038
          36921 => x"80", -- $09039
          36922 => x"80", -- $0903a
          36923 => x"80", -- $0903b
          36924 => x"80", -- $0903c
          36925 => x"80", -- $0903d
          36926 => x"80", -- $0903e
          36927 => x"80", -- $0903f
          36928 => x"80", -- $09040
          36929 => x"80", -- $09041
          36930 => x"80", -- $09042
          36931 => x"81", -- $09043
          36932 => x"80", -- $09044
          36933 => x"80", -- $09045
          36934 => x"80", -- $09046
          36935 => x"80", -- $09047
          36936 => x"80", -- $09048
          36937 => x"80", -- $09049
          36938 => x"80", -- $0904a
          36939 => x"80", -- $0904b
          36940 => x"80", -- $0904c
          36941 => x"80", -- $0904d
          36942 => x"80", -- $0904e
          36943 => x"80", -- $0904f
          36944 => x"80", -- $09050
          36945 => x"80", -- $09051
          36946 => x"80", -- $09052
          36947 => x"80", -- $09053
          36948 => x"80", -- $09054
          36949 => x"80", -- $09055
          36950 => x"80", -- $09056
          36951 => x"80", -- $09057
          36952 => x"80", -- $09058
          36953 => x"80", -- $09059
          36954 => x"80", -- $0905a
          36955 => x"80", -- $0905b
          36956 => x"80", -- $0905c
          36957 => x"80", -- $0905d
          36958 => x"80", -- $0905e
          36959 => x"80", -- $0905f
          36960 => x"80", -- $09060
          36961 => x"80", -- $09061
          36962 => x"80", -- $09062
          36963 => x"80", -- $09063
          36964 => x"80", -- $09064
          36965 => x"80", -- $09065
          36966 => x"80", -- $09066
          36967 => x"80", -- $09067
          36968 => x"80", -- $09068
          36969 => x"80", -- $09069
          36970 => x"80", -- $0906a
          36971 => x"80", -- $0906b
          36972 => x"80", -- $0906c
          36973 => x"80", -- $0906d
          36974 => x"80", -- $0906e
          36975 => x"80", -- $0906f
          36976 => x"80", -- $09070
          36977 => x"80", -- $09071
          36978 => x"80", -- $09072
          36979 => x"80", -- $09073
          36980 => x"80", -- $09074
          36981 => x"80", -- $09075
          36982 => x"80", -- $09076
          36983 => x"80", -- $09077
          36984 => x"80", -- $09078
          36985 => x"80", -- $09079
          36986 => x"80", -- $0907a
          36987 => x"80", -- $0907b
          36988 => x"80", -- $0907c
          36989 => x"80", -- $0907d
          36990 => x"80", -- $0907e
          36991 => x"80", -- $0907f
          36992 => x"80", -- $09080
          36993 => x"80", -- $09081
          36994 => x"80", -- $09082
          36995 => x"80", -- $09083
          36996 => x"80", -- $09084
          36997 => x"80", -- $09085
          36998 => x"80", -- $09086
          36999 => x"80", -- $09087
          37000 => x"80", -- $09088
          37001 => x"80", -- $09089
          37002 => x"80", -- $0908a
          37003 => x"80", -- $0908b
          37004 => x"80", -- $0908c
          37005 => x"80", -- $0908d
          37006 => x"80", -- $0908e
          37007 => x"80", -- $0908f
          37008 => x"80", -- $09090
          37009 => x"80", -- $09091
          37010 => x"80", -- $09092
          37011 => x"80", -- $09093
          37012 => x"80", -- $09094
          37013 => x"80", -- $09095
          37014 => x"80", -- $09096
          37015 => x"80", -- $09097
          37016 => x"80", -- $09098
          37017 => x"80", -- $09099
          37018 => x"80", -- $0909a
          37019 => x"80", -- $0909b
          37020 => x"80", -- $0909c
          37021 => x"80", -- $0909d
          37022 => x"80", -- $0909e
          37023 => x"80", -- $0909f
          37024 => x"80", -- $090a0
          37025 => x"80", -- $090a1
          37026 => x"80", -- $090a2
          37027 => x"80", -- $090a3
          37028 => x"80", -- $090a4
          37029 => x"80", -- $090a5
          37030 => x"80", -- $090a6
          37031 => x"80", -- $090a7
          37032 => x"80", -- $090a8
          37033 => x"80", -- $090a9
          37034 => x"80", -- $090aa
          37035 => x"80", -- $090ab
          37036 => x"80", -- $090ac
          37037 => x"80", -- $090ad
          37038 => x"80", -- $090ae
          37039 => x"80", -- $090af
          37040 => x"80", -- $090b0
          37041 => x"80", -- $090b1
          37042 => x"80", -- $090b2
          37043 => x"80", -- $090b3
          37044 => x"80", -- $090b4
          37045 => x"80", -- $090b5
          37046 => x"80", -- $090b6
          37047 => x"80", -- $090b7
          37048 => x"80", -- $090b8
          37049 => x"80", -- $090b9
          37050 => x"80", -- $090ba
          37051 => x"80", -- $090bb
          37052 => x"80", -- $090bc
          37053 => x"80", -- $090bd
          37054 => x"80", -- $090be
          37055 => x"80", -- $090bf
          37056 => x"80", -- $090c0
          37057 => x"80", -- $090c1
          37058 => x"80", -- $090c2
          37059 => x"80", -- $090c3
          37060 => x"80", -- $090c4
          37061 => x"80", -- $090c5
          37062 => x"80", -- $090c6
          37063 => x"80", -- $090c7
          37064 => x"80", -- $090c8
          37065 => x"80", -- $090c9
          37066 => x"80", -- $090ca
          37067 => x"80", -- $090cb
          37068 => x"80", -- $090cc
          37069 => x"80", -- $090cd
          37070 => x"80", -- $090ce
          37071 => x"80", -- $090cf
          37072 => x"80", -- $090d0
          37073 => x"80", -- $090d1
          37074 => x"80", -- $090d2
          37075 => x"80", -- $090d3
          37076 => x"80", -- $090d4
          37077 => x"80", -- $090d5
          37078 => x"80", -- $090d6
          37079 => x"80", -- $090d7
          37080 => x"80", -- $090d8
          37081 => x"80", -- $090d9
          37082 => x"80", -- $090da
          37083 => x"80", -- $090db
          37084 => x"80", -- $090dc
          37085 => x"80", -- $090dd
          37086 => x"80", -- $090de
          37087 => x"80", -- $090df
          37088 => x"80", -- $090e0
          37089 => x"80", -- $090e1
          37090 => x"80", -- $090e2
          37091 => x"80", -- $090e3
          37092 => x"80", -- $090e4
          37093 => x"80", -- $090e5
          37094 => x"80", -- $090e6
          37095 => x"80", -- $090e7
          37096 => x"80", -- $090e8
          37097 => x"80", -- $090e9
          37098 => x"80", -- $090ea
          37099 => x"80", -- $090eb
          37100 => x"80", -- $090ec
          37101 => x"80", -- $090ed
          37102 => x"80", -- $090ee
          37103 => x"80", -- $090ef
          37104 => x"80", -- $090f0
          37105 => x"80", -- $090f1
          37106 => x"80", -- $090f2
          37107 => x"80", -- $090f3
          37108 => x"80", -- $090f4
          37109 => x"80", -- $090f5
          37110 => x"80", -- $090f6
          37111 => x"80", -- $090f7
          37112 => x"80", -- $090f8
          37113 => x"80", -- $090f9
          37114 => x"80", -- $090fa
          37115 => x"80", -- $090fb
          37116 => x"80", -- $090fc
          37117 => x"80", -- $090fd
          37118 => x"80", -- $090fe
          37119 => x"80", -- $090ff
          37120 => x"80", -- $09100
          37121 => x"80", -- $09101
          37122 => x"80", -- $09102
          37123 => x"80", -- $09103
          37124 => x"80", -- $09104
          37125 => x"80", -- $09105
          37126 => x"80", -- $09106
          37127 => x"80", -- $09107
          37128 => x"80", -- $09108
          37129 => x"80", -- $09109
          37130 => x"80", -- $0910a
          37131 => x"80", -- $0910b
          37132 => x"80", -- $0910c
          37133 => x"80", -- $0910d
          37134 => x"80", -- $0910e
          37135 => x"80", -- $0910f
          37136 => x"80", -- $09110
          37137 => x"80", -- $09111
          37138 => x"80", -- $09112
          37139 => x"80", -- $09113
          37140 => x"80", -- $09114
          37141 => x"80", -- $09115
          37142 => x"80", -- $09116
          37143 => x"80", -- $09117
          37144 => x"80", -- $09118
          37145 => x"80", -- $09119
          37146 => x"80", -- $0911a
          37147 => x"80", -- $0911b
          37148 => x"80", -- $0911c
          37149 => x"80", -- $0911d
          37150 => x"80", -- $0911e
          37151 => x"80", -- $0911f
          37152 => x"80", -- $09120
          37153 => x"80", -- $09121
          37154 => x"80", -- $09122
          37155 => x"80", -- $09123
          37156 => x"80", -- $09124
          37157 => x"80", -- $09125
          37158 => x"80", -- $09126
          37159 => x"80", -- $09127
          37160 => x"80", -- $09128
          37161 => x"80", -- $09129
          37162 => x"80", -- $0912a
          37163 => x"80", -- $0912b
          37164 => x"80", -- $0912c
          37165 => x"80", -- $0912d
          37166 => x"80", -- $0912e
          37167 => x"80", -- $0912f
          37168 => x"80", -- $09130
          37169 => x"80", -- $09131
          37170 => x"80", -- $09132
          37171 => x"80", -- $09133
          37172 => x"80", -- $09134
          37173 => x"80", -- $09135
          37174 => x"80", -- $09136
          37175 => x"80", -- $09137
          37176 => x"80", -- $09138
          37177 => x"80", -- $09139
          37178 => x"80", -- $0913a
          37179 => x"80", -- $0913b
          37180 => x"80", -- $0913c
          37181 => x"80", -- $0913d
          37182 => x"80", -- $0913e
          37183 => x"80", -- $0913f
          37184 => x"80", -- $09140
          37185 => x"80", -- $09141
          37186 => x"80", -- $09142
          37187 => x"80", -- $09143
          37188 => x"80", -- $09144
          37189 => x"80", -- $09145
          37190 => x"80", -- $09146
          37191 => x"80", -- $09147
          37192 => x"80", -- $09148
          37193 => x"80", -- $09149
          37194 => x"80", -- $0914a
          37195 => x"80", -- $0914b
          37196 => x"80", -- $0914c
          37197 => x"80", -- $0914d
          37198 => x"80", -- $0914e
          37199 => x"80", -- $0914f
          37200 => x"80", -- $09150
          37201 => x"80", -- $09151
          37202 => x"80", -- $09152
          37203 => x"80", -- $09153
          37204 => x"80", -- $09154
          37205 => x"80", -- $09155
          37206 => x"80", -- $09156
          37207 => x"80", -- $09157
          37208 => x"80", -- $09158
          37209 => x"7f", -- $09159
          37210 => x"7f", -- $0915a
          37211 => x"7f", -- $0915b
          37212 => x"7f", -- $0915c
          37213 => x"7f", -- $0915d
          37214 => x"7f", -- $0915e
          37215 => x"7f", -- $0915f
          37216 => x"7f", -- $09160
          37217 => x"7f", -- $09161
          37218 => x"7f", -- $09162
          37219 => x"7f", -- $09163
          37220 => x"80", -- $09164
          37221 => x"80", -- $09165
          37222 => x"80", -- $09166
          37223 => x"80", -- $09167
          37224 => x"80", -- $09168
          37225 => x"80", -- $09169
          37226 => x"80", -- $0916a
          37227 => x"80", -- $0916b
          37228 => x"80", -- $0916c
          37229 => x"80", -- $0916d
          37230 => x"80", -- $0916e
          37231 => x"80", -- $0916f
          37232 => x"80", -- $09170
          37233 => x"80", -- $09171
          37234 => x"80", -- $09172
          37235 => x"80", -- $09173
          37236 => x"7f", -- $09174
          37237 => x"80", -- $09175
          37238 => x"7f", -- $09176
          37239 => x"7f", -- $09177
          37240 => x"7f", -- $09178
          37241 => x"7f", -- $09179
          37242 => x"7f", -- $0917a
          37243 => x"7f", -- $0917b
          37244 => x"7f", -- $0917c
          37245 => x"7f", -- $0917d
          37246 => x"7f", -- $0917e
          37247 => x"7f", -- $0917f
          37248 => x"7f", -- $09180
          37249 => x"7f", -- $09181
          37250 => x"7f", -- $09182
          37251 => x"7f", -- $09183
          37252 => x"80", -- $09184
          37253 => x"80", -- $09185
          37254 => x"80", -- $09186
          37255 => x"80", -- $09187
          37256 => x"80", -- $09188
          37257 => x"80", -- $09189
          37258 => x"80", -- $0918a
          37259 => x"80", -- $0918b
          37260 => x"80", -- $0918c
          37261 => x"80", -- $0918d
          37262 => x"80", -- $0918e
          37263 => x"80", -- $0918f
          37264 => x"80", -- $09190
          37265 => x"80", -- $09191
          37266 => x"80", -- $09192
          37267 => x"80", -- $09193
          37268 => x"80", -- $09194
          37269 => x"80", -- $09195
          37270 => x"80", -- $09196
          37271 => x"80", -- $09197
          37272 => x"80", -- $09198
          37273 => x"80", -- $09199
          37274 => x"80", -- $0919a
          37275 => x"7f", -- $0919b
          37276 => x"7f", -- $0919c
          37277 => x"7f", -- $0919d
          37278 => x"7f", -- $0919e
          37279 => x"7f", -- $0919f
          37280 => x"7f", -- $091a0
          37281 => x"80", -- $091a1
          37282 => x"80", -- $091a2
          37283 => x"80", -- $091a3
          37284 => x"80", -- $091a4
          37285 => x"80", -- $091a5
          37286 => x"80", -- $091a6
          37287 => x"80", -- $091a7
          37288 => x"80", -- $091a8
          37289 => x"80", -- $091a9
          37290 => x"80", -- $091aa
          37291 => x"80", -- $091ab
          37292 => x"80", -- $091ac
          37293 => x"80", -- $091ad
          37294 => x"80", -- $091ae
          37295 => x"80", -- $091af
          37296 => x"80", -- $091b0
          37297 => x"80", -- $091b1
          37298 => x"80", -- $091b2
          37299 => x"80", -- $091b3
          37300 => x"80", -- $091b4
          37301 => x"80", -- $091b5
          37302 => x"80", -- $091b6
          37303 => x"80", -- $091b7
          37304 => x"80", -- $091b8
          37305 => x"80", -- $091b9
          37306 => x"80", -- $091ba
          37307 => x"80", -- $091bb
          37308 => x"80", -- $091bc
          37309 => x"80", -- $091bd
          37310 => x"80", -- $091be
          37311 => x"80", -- $091bf
          37312 => x"80", -- $091c0
          37313 => x"80", -- $091c1
          37314 => x"80", -- $091c2
          37315 => x"80", -- $091c3
          37316 => x"80", -- $091c4
          37317 => x"80", -- $091c5
          37318 => x"80", -- $091c6
          37319 => x"80", -- $091c7
          37320 => x"80", -- $091c8
          37321 => x"80", -- $091c9
          37322 => x"80", -- $091ca
          37323 => x"80", -- $091cb
          37324 => x"80", -- $091cc
          37325 => x"80", -- $091cd
          37326 => x"80", -- $091ce
          37327 => x"80", -- $091cf
          37328 => x"80", -- $091d0
          37329 => x"80", -- $091d1
          37330 => x"80", -- $091d2
          37331 => x"80", -- $091d3
          37332 => x"80", -- $091d4
          37333 => x"80", -- $091d5
          37334 => x"80", -- $091d6
          37335 => x"80", -- $091d7
          37336 => x"80", -- $091d8
          37337 => x"80", -- $091d9
          37338 => x"80", -- $091da
          37339 => x"80", -- $091db
          37340 => x"80", -- $091dc
          37341 => x"80", -- $091dd
          37342 => x"80", -- $091de
          37343 => x"80", -- $091df
          37344 => x"80", -- $091e0
          37345 => x"80", -- $091e1
          37346 => x"80", -- $091e2
          37347 => x"80", -- $091e3
          37348 => x"80", -- $091e4
          37349 => x"80", -- $091e5
          37350 => x"80", -- $091e6
          37351 => x"80", -- $091e7
          37352 => x"80", -- $091e8
          37353 => x"80", -- $091e9
          37354 => x"80", -- $091ea
          37355 => x"80", -- $091eb
          37356 => x"81", -- $091ec
          37357 => x"81", -- $091ed
          37358 => x"80", -- $091ee
          37359 => x"81", -- $091ef
          37360 => x"81", -- $091f0
          37361 => x"80", -- $091f1
          37362 => x"80", -- $091f2
          37363 => x"80", -- $091f3
          37364 => x"80", -- $091f4
          37365 => x"80", -- $091f5
          37366 => x"80", -- $091f6
          37367 => x"80", -- $091f7
          37368 => x"80", -- $091f8
          37369 => x"80", -- $091f9
          37370 => x"80", -- $091fa
          37371 => x"80", -- $091fb
          37372 => x"80", -- $091fc
          37373 => x"80", -- $091fd
          37374 => x"80", -- $091fe
          37375 => x"80", -- $091ff
          37376 => x"80", -- $09200
          37377 => x"80", -- $09201
          37378 => x"80", -- $09202
          37379 => x"80", -- $09203
          37380 => x"80", -- $09204
          37381 => x"80", -- $09205
          37382 => x"80", -- $09206
          37383 => x"80", -- $09207
          37384 => x"80", -- $09208
          37385 => x"80", -- $09209
          37386 => x"80", -- $0920a
          37387 => x"80", -- $0920b
          37388 => x"80", -- $0920c
          37389 => x"80", -- $0920d
          37390 => x"80", -- $0920e
          37391 => x"80", -- $0920f
          37392 => x"80", -- $09210
          37393 => x"80", -- $09211
          37394 => x"80", -- $09212
          37395 => x"80", -- $09213
          37396 => x"80", -- $09214
          37397 => x"80", -- $09215
          37398 => x"80", -- $09216
          37399 => x"80", -- $09217
          37400 => x"80", -- $09218
          37401 => x"80", -- $09219
          37402 => x"80", -- $0921a
          37403 => x"80", -- $0921b
          37404 => x"80", -- $0921c
          37405 => x"80", -- $0921d
          37406 => x"80", -- $0921e
          37407 => x"80", -- $0921f
          37408 => x"80", -- $09220
          37409 => x"80", -- $09221
          37410 => x"80", -- $09222
          37411 => x"80", -- $09223
          37412 => x"80", -- $09224
          37413 => x"80", -- $09225
          37414 => x"80", -- $09226
          37415 => x"80", -- $09227
          37416 => x"80", -- $09228
          37417 => x"80", -- $09229
          37418 => x"80", -- $0922a
          37419 => x"80", -- $0922b
          37420 => x"80", -- $0922c
          37421 => x"80", -- $0922d
          37422 => x"80", -- $0922e
          37423 => x"80", -- $0922f
          37424 => x"80", -- $09230
          37425 => x"80", -- $09231
          37426 => x"80", -- $09232
          37427 => x"80", -- $09233
          37428 => x"80", -- $09234
          37429 => x"80", -- $09235
          37430 => x"80", -- $09236
          37431 => x"80", -- $09237
          37432 => x"80", -- $09238
          37433 => x"80", -- $09239
          37434 => x"80", -- $0923a
          37435 => x"80", -- $0923b
          37436 => x"80", -- $0923c
          37437 => x"80", -- $0923d
          37438 => x"80", -- $0923e
          37439 => x"80", -- $0923f
          37440 => x"80", -- $09240
          37441 => x"80", -- $09241
          37442 => x"80", -- $09242
          37443 => x"80", -- $09243
          37444 => x"80", -- $09244
          37445 => x"80", -- $09245
          37446 => x"80", -- $09246
          37447 => x"80", -- $09247
          37448 => x"80", -- $09248
          37449 => x"80", -- $09249
          37450 => x"80", -- $0924a
          37451 => x"80", -- $0924b
          37452 => x"80", -- $0924c
          37453 => x"80", -- $0924d
          37454 => x"80", -- $0924e
          37455 => x"80", -- $0924f
          37456 => x"80", -- $09250
          37457 => x"80", -- $09251
          37458 => x"80", -- $09252
          37459 => x"80", -- $09253
          37460 => x"80", -- $09254
          37461 => x"80", -- $09255
          37462 => x"80", -- $09256
          37463 => x"80", -- $09257
          37464 => x"80", -- $09258
          37465 => x"80", -- $09259
          37466 => x"80", -- $0925a
          37467 => x"80", -- $0925b
          37468 => x"80", -- $0925c
          37469 => x"80", -- $0925d
          37470 => x"80", -- $0925e
          37471 => x"80", -- $0925f
          37472 => x"80", -- $09260
          37473 => x"80", -- $09261
          37474 => x"80", -- $09262
          37475 => x"80", -- $09263
          37476 => x"80", -- $09264
          37477 => x"80", -- $09265
          37478 => x"80", -- $09266
          37479 => x"80", -- $09267
          37480 => x"80", -- $09268
          37481 => x"80", -- $09269
          37482 => x"80", -- $0926a
          37483 => x"80", -- $0926b
          37484 => x"80", -- $0926c
          37485 => x"80", -- $0926d
          37486 => x"80", -- $0926e
          37487 => x"80", -- $0926f
          37488 => x"80", -- $09270
          37489 => x"80", -- $09271
          37490 => x"80", -- $09272
          37491 => x"80", -- $09273
          37492 => x"80", -- $09274
          37493 => x"80", -- $09275
          37494 => x"80", -- $09276
          37495 => x"80", -- $09277
          37496 => x"80", -- $09278
          37497 => x"80", -- $09279
          37498 => x"80", -- $0927a
          37499 => x"80", -- $0927b
          37500 => x"80", -- $0927c
          37501 => x"80", -- $0927d
          37502 => x"80", -- $0927e
          37503 => x"80", -- $0927f
          37504 => x"80", -- $09280
          37505 => x"80", -- $09281
          37506 => x"80", -- $09282
          37507 => x"80", -- $09283
          37508 => x"80", -- $09284
          37509 => x"80", -- $09285
          37510 => x"80", -- $09286
          37511 => x"80", -- $09287
          37512 => x"80", -- $09288
          37513 => x"80", -- $09289
          37514 => x"80", -- $0928a
          37515 => x"80", -- $0928b
          37516 => x"80", -- $0928c
          37517 => x"80", -- $0928d
          37518 => x"80", -- $0928e
          37519 => x"80", -- $0928f
          37520 => x"80", -- $09290
          37521 => x"80", -- $09291
          37522 => x"80", -- $09292
          37523 => x"80", -- $09293
          37524 => x"80", -- $09294
          37525 => x"80", -- $09295
          37526 => x"80", -- $09296
          37527 => x"80", -- $09297
          37528 => x"80", -- $09298
          37529 => x"80", -- $09299
          37530 => x"80", -- $0929a
          37531 => x"80", -- $0929b
          37532 => x"80", -- $0929c
          37533 => x"80", -- $0929d
          37534 => x"80", -- $0929e
          37535 => x"80", -- $0929f
          37536 => x"80", -- $092a0
          37537 => x"80", -- $092a1
          37538 => x"80", -- $092a2
          37539 => x"80", -- $092a3
          37540 => x"80", -- $092a4
          37541 => x"80", -- $092a5
          37542 => x"80", -- $092a6
          37543 => x"80", -- $092a7
          37544 => x"80", -- $092a8
          37545 => x"80", -- $092a9
          37546 => x"80", -- $092aa
          37547 => x"81", -- $092ab
          37548 => x"81", -- $092ac
          37549 => x"81", -- $092ad
          37550 => x"81", -- $092ae
          37551 => x"81", -- $092af
          37552 => x"81", -- $092b0
          37553 => x"81", -- $092b1
          37554 => x"81", -- $092b2
          37555 => x"81", -- $092b3
          37556 => x"80", -- $092b4
          37557 => x"80", -- $092b5
          37558 => x"80", -- $092b6
          37559 => x"80", -- $092b7
          37560 => x"80", -- $092b8
          37561 => x"80", -- $092b9
          37562 => x"80", -- $092ba
          37563 => x"80", -- $092bb
          37564 => x"80", -- $092bc
          37565 => x"80", -- $092bd
          37566 => x"80", -- $092be
          37567 => x"80", -- $092bf
          37568 => x"80", -- $092c0
          37569 => x"80", -- $092c1
          37570 => x"81", -- $092c2
          37571 => x"81", -- $092c3
          37572 => x"81", -- $092c4
          37573 => x"81", -- $092c5
          37574 => x"81", -- $092c6
          37575 => x"81", -- $092c7
          37576 => x"81", -- $092c8
          37577 => x"81", -- $092c9
          37578 => x"81", -- $092ca
          37579 => x"81", -- $092cb
          37580 => x"81", -- $092cc
          37581 => x"81", -- $092cd
          37582 => x"81", -- $092ce
          37583 => x"81", -- $092cf
          37584 => x"81", -- $092d0
          37585 => x"81", -- $092d1
          37586 => x"81", -- $092d2
          37587 => x"81", -- $092d3
          37588 => x"81", -- $092d4
          37589 => x"81", -- $092d5
          37590 => x"81", -- $092d6
          37591 => x"80", -- $092d7
          37592 => x"80", -- $092d8
          37593 => x"80", -- $092d9
          37594 => x"80", -- $092da
          37595 => x"80", -- $092db
          37596 => x"80", -- $092dc
          37597 => x"80", -- $092dd
          37598 => x"80", -- $092de
          37599 => x"80", -- $092df
          37600 => x"80", -- $092e0
          37601 => x"80", -- $092e1
          37602 => x"80", -- $092e2
          37603 => x"80", -- $092e3
          37604 => x"80", -- $092e4
          37605 => x"81", -- $092e5
          37606 => x"81", -- $092e6
          37607 => x"81", -- $092e7
          37608 => x"81", -- $092e8
          37609 => x"81", -- $092e9
          37610 => x"81", -- $092ea
          37611 => x"81", -- $092eb
          37612 => x"81", -- $092ec
          37613 => x"81", -- $092ed
          37614 => x"81", -- $092ee
          37615 => x"81", -- $092ef
          37616 => x"81", -- $092f0
          37617 => x"81", -- $092f1
          37618 => x"81", -- $092f2
          37619 => x"81", -- $092f3
          37620 => x"81", -- $092f4
          37621 => x"80", -- $092f5
          37622 => x"80", -- $092f6
          37623 => x"80", -- $092f7
          37624 => x"80", -- $092f8
          37625 => x"80", -- $092f9
          37626 => x"80", -- $092fa
          37627 => x"80", -- $092fb
          37628 => x"80", -- $092fc
          37629 => x"80", -- $092fd
          37630 => x"80", -- $092fe
          37631 => x"80", -- $092ff
          37632 => x"80", -- $09300
          37633 => x"80", -- $09301
          37634 => x"80", -- $09302
          37635 => x"80", -- $09303
          37636 => x"80", -- $09304
          37637 => x"81", -- $09305
          37638 => x"81", -- $09306
          37639 => x"80", -- $09307
          37640 => x"80", -- $09308
          37641 => x"80", -- $09309
          37642 => x"80", -- $0930a
          37643 => x"80", -- $0930b
          37644 => x"80", -- $0930c
          37645 => x"80", -- $0930d
          37646 => x"80", -- $0930e
          37647 => x"80", -- $0930f
          37648 => x"80", -- $09310
          37649 => x"80", -- $09311
          37650 => x"80", -- $09312
          37651 => x"80", -- $09313
          37652 => x"80", -- $09314
          37653 => x"80", -- $09315
          37654 => x"80", -- $09316
          37655 => x"80", -- $09317
          37656 => x"80", -- $09318
          37657 => x"80", -- $09319
          37658 => x"80", -- $0931a
          37659 => x"80", -- $0931b
          37660 => x"80", -- $0931c
          37661 => x"80", -- $0931d
          37662 => x"80", -- $0931e
          37663 => x"80", -- $0931f
          37664 => x"80", -- $09320
          37665 => x"80", -- $09321
          37666 => x"80", -- $09322
          37667 => x"80", -- $09323
          37668 => x"80", -- $09324
          37669 => x"80", -- $09325
          37670 => x"80", -- $09326
          37671 => x"80", -- $09327
          37672 => x"80", -- $09328
          37673 => x"80", -- $09329
          37674 => x"80", -- $0932a
          37675 => x"80", -- $0932b
          37676 => x"80", -- $0932c
          37677 => x"80", -- $0932d
          37678 => x"80", -- $0932e
          37679 => x"80", -- $0932f
          37680 => x"80", -- $09330
          37681 => x"80", -- $09331
          37682 => x"80", -- $09332
          37683 => x"80", -- $09333
          37684 => x"80", -- $09334
          37685 => x"80", -- $09335
          37686 => x"80", -- $09336
          37687 => x"80", -- $09337
          37688 => x"80", -- $09338
          37689 => x"80", -- $09339
          37690 => x"80", -- $0933a
          37691 => x"80", -- $0933b
          37692 => x"80", -- $0933c
          37693 => x"80", -- $0933d
          37694 => x"80", -- $0933e
          37695 => x"80", -- $0933f
          37696 => x"80", -- $09340
          37697 => x"80", -- $09341
          37698 => x"80", -- $09342
          37699 => x"80", -- $09343
          37700 => x"80", -- $09344
          37701 => x"80", -- $09345
          37702 => x"80", -- $09346
          37703 => x"80", -- $09347
          37704 => x"80", -- $09348
          37705 => x"80", -- $09349
          37706 => x"80", -- $0934a
          37707 => x"80", -- $0934b
          37708 => x"80", -- $0934c
          37709 => x"80", -- $0934d
          37710 => x"80", -- $0934e
          37711 => x"80", -- $0934f
          37712 => x"80", -- $09350
          37713 => x"80", -- $09351
          37714 => x"80", -- $09352
          37715 => x"80", -- $09353
          37716 => x"80", -- $09354
          37717 => x"80", -- $09355
          37718 => x"7f", -- $09356
          37719 => x"7f", -- $09357
          37720 => x"7f", -- $09358
          37721 => x"7f", -- $09359
          37722 => x"80", -- $0935a
          37723 => x"80", -- $0935b
          37724 => x"80", -- $0935c
          37725 => x"80", -- $0935d
          37726 => x"80", -- $0935e
          37727 => x"80", -- $0935f
          37728 => x"80", -- $09360
          37729 => x"80", -- $09361
          37730 => x"80", -- $09362
          37731 => x"80", -- $09363
          37732 => x"80", -- $09364
          37733 => x"80", -- $09365
          37734 => x"80", -- $09366
          37735 => x"80", -- $09367
          37736 => x"80", -- $09368
          37737 => x"80", -- $09369
          37738 => x"80", -- $0936a
          37739 => x"80", -- $0936b
          37740 => x"80", -- $0936c
          37741 => x"80", -- $0936d
          37742 => x"80", -- $0936e
          37743 => x"80", -- $0936f
          37744 => x"80", -- $09370
          37745 => x"80", -- $09371
          37746 => x"80", -- $09372
          37747 => x"80", -- $09373
          37748 => x"80", -- $09374
          37749 => x"80", -- $09375
          37750 => x"80", -- $09376
          37751 => x"80", -- $09377
          37752 => x"80", -- $09378
          37753 => x"80", -- $09379
          37754 => x"80", -- $0937a
          37755 => x"80", -- $0937b
          37756 => x"80", -- $0937c
          37757 => x"80", -- $0937d
          37758 => x"80", -- $0937e
          37759 => x"80", -- $0937f
          37760 => x"80", -- $09380
          37761 => x"80", -- $09381
          37762 => x"80", -- $09382
          37763 => x"80", -- $09383
          37764 => x"80", -- $09384
          37765 => x"80", -- $09385
          37766 => x"80", -- $09386
          37767 => x"80", -- $09387
          37768 => x"80", -- $09388
          37769 => x"80", -- $09389
          37770 => x"80", -- $0938a
          37771 => x"80", -- $0938b
          37772 => x"80", -- $0938c
          37773 => x"80", -- $0938d
          37774 => x"80", -- $0938e
          37775 => x"80", -- $0938f
          37776 => x"80", -- $09390
          37777 => x"80", -- $09391
          37778 => x"80", -- $09392
          37779 => x"80", -- $09393
          37780 => x"80", -- $09394
          37781 => x"80", -- $09395
          37782 => x"80", -- $09396
          37783 => x"80", -- $09397
          37784 => x"80", -- $09398
          37785 => x"80", -- $09399
          37786 => x"80", -- $0939a
          37787 => x"80", -- $0939b
          37788 => x"80", -- $0939c
          37789 => x"80", -- $0939d
          37790 => x"80", -- $0939e
          37791 => x"80", -- $0939f
          37792 => x"80", -- $093a0
          37793 => x"80", -- $093a1
          37794 => x"80", -- $093a2
          37795 => x"80", -- $093a3
          37796 => x"80", -- $093a4
          37797 => x"80", -- $093a5
          37798 => x"80", -- $093a6
          37799 => x"80", -- $093a7
          37800 => x"80", -- $093a8
          37801 => x"80", -- $093a9
          37802 => x"80", -- $093aa
          37803 => x"80", -- $093ab
          37804 => x"80", -- $093ac
          37805 => x"80", -- $093ad
          37806 => x"80", -- $093ae
          37807 => x"80", -- $093af
          37808 => x"80", -- $093b0
          37809 => x"80", -- $093b1
          37810 => x"80", -- $093b2
          37811 => x"80", -- $093b3
          37812 => x"80", -- $093b4
          37813 => x"80", -- $093b5
          37814 => x"80", -- $093b6
          37815 => x"80", -- $093b7
          37816 => x"80", -- $093b8
          37817 => x"80", -- $093b9
          37818 => x"80", -- $093ba
          37819 => x"80", -- $093bb
          37820 => x"80", -- $093bc
          37821 => x"80", -- $093bd
          37822 => x"80", -- $093be
          37823 => x"80", -- $093bf
          37824 => x"80", -- $093c0
          37825 => x"80", -- $093c1
          37826 => x"80", -- $093c2
          37827 => x"80", -- $093c3
          37828 => x"80", -- $093c4
          37829 => x"80", -- $093c5
          37830 => x"80", -- $093c6
          37831 => x"80", -- $093c7
          37832 => x"80", -- $093c8
          37833 => x"80", -- $093c9
          37834 => x"80", -- $093ca
          37835 => x"80", -- $093cb
          37836 => x"80", -- $093cc
          37837 => x"80", -- $093cd
          37838 => x"80", -- $093ce
          37839 => x"80", -- $093cf
          37840 => x"80", -- $093d0
          37841 => x"80", -- $093d1
          37842 => x"80", -- $093d2
          37843 => x"80", -- $093d3
          37844 => x"80", -- $093d4
          37845 => x"80", -- $093d5
          37846 => x"80", -- $093d6
          37847 => x"80", -- $093d7
          37848 => x"80", -- $093d8
          37849 => x"80", -- $093d9
          37850 => x"80", -- $093da
          37851 => x"80", -- $093db
          37852 => x"7f", -- $093dc
          37853 => x"80", -- $093dd
          37854 => x"80", -- $093de
          37855 => x"80", -- $093df
          37856 => x"80", -- $093e0
          37857 => x"80", -- $093e1
          37858 => x"7f", -- $093e2
          37859 => x"7f", -- $093e3
          37860 => x"7f", -- $093e4
          37861 => x"7f", -- $093e5
          37862 => x"7f", -- $093e6
          37863 => x"7f", -- $093e7
          37864 => x"7f", -- $093e8
          37865 => x"7f", -- $093e9
          37866 => x"7f", -- $093ea
          37867 => x"7f", -- $093eb
          37868 => x"7f", -- $093ec
          37869 => x"7f", -- $093ed
          37870 => x"80", -- $093ee
          37871 => x"7f", -- $093ef
          37872 => x"7f", -- $093f0
          37873 => x"7f", -- $093f1
          37874 => x"7f", -- $093f2
          37875 => x"7f", -- $093f3
          37876 => x"7f", -- $093f4
          37877 => x"7f", -- $093f5
          37878 => x"7f", -- $093f6
          37879 => x"80", -- $093f7
          37880 => x"80", -- $093f8
          37881 => x"80", -- $093f9
          37882 => x"80", -- $093fa
          37883 => x"80", -- $093fb
          37884 => x"80", -- $093fc
          37885 => x"80", -- $093fd
          37886 => x"80", -- $093fe
          37887 => x"80", -- $093ff
          37888 => x"80", -- $09400
          37889 => x"80", -- $09401
          37890 => x"80", -- $09402
          37891 => x"7f", -- $09403
          37892 => x"7f", -- $09404
          37893 => x"7f", -- $09405
          37894 => x"7f", -- $09406
          37895 => x"80", -- $09407
          37896 => x"80", -- $09408
          37897 => x"80", -- $09409
          37898 => x"80", -- $0940a
          37899 => x"80", -- $0940b
          37900 => x"80", -- $0940c
          37901 => x"80", -- $0940d
          37902 => x"80", -- $0940e
          37903 => x"80", -- $0940f
          37904 => x"80", -- $09410
          37905 => x"80", -- $09411
          37906 => x"80", -- $09412
          37907 => x"80", -- $09413
          37908 => x"80", -- $09414
          37909 => x"80", -- $09415
          37910 => x"80", -- $09416
          37911 => x"80", -- $09417
          37912 => x"80", -- $09418
          37913 => x"80", -- $09419
          37914 => x"80", -- $0941a
          37915 => x"80", -- $0941b
          37916 => x"80", -- $0941c
          37917 => x"80", -- $0941d
          37918 => x"80", -- $0941e
          37919 => x"80", -- $0941f
          37920 => x"80", -- $09420
          37921 => x"80", -- $09421
          37922 => x"80", -- $09422
          37923 => x"80", -- $09423
          37924 => x"80", -- $09424
          37925 => x"80", -- $09425
          37926 => x"80", -- $09426
          37927 => x"80", -- $09427
          37928 => x"80", -- $09428
          37929 => x"80", -- $09429
          37930 => x"80", -- $0942a
          37931 => x"80", -- $0942b
          37932 => x"80", -- $0942c
          37933 => x"80", -- $0942d
          37934 => x"80", -- $0942e
          37935 => x"80", -- $0942f
          37936 => x"80", -- $09430
          37937 => x"80", -- $09431
          37938 => x"80", -- $09432
          37939 => x"80", -- $09433
          37940 => x"80", -- $09434
          37941 => x"80", -- $09435
          37942 => x"80", -- $09436
          37943 => x"80", -- $09437
          37944 => x"80", -- $09438
          37945 => x"80", -- $09439
          37946 => x"80", -- $0943a
          37947 => x"80", -- $0943b
          37948 => x"80", -- $0943c
          37949 => x"80", -- $0943d
          37950 => x"80", -- $0943e
          37951 => x"80", -- $0943f
          37952 => x"80", -- $09440
          37953 => x"80", -- $09441
          37954 => x"80", -- $09442
          37955 => x"80", -- $09443
          37956 => x"80", -- $09444
          37957 => x"80", -- $09445
          37958 => x"80", -- $09446
          37959 => x"80", -- $09447
          37960 => x"80", -- $09448
          37961 => x"80", -- $09449
          37962 => x"80", -- $0944a
          37963 => x"80", -- $0944b
          37964 => x"80", -- $0944c
          37965 => x"80", -- $0944d
          37966 => x"80", -- $0944e
          37967 => x"80", -- $0944f
          37968 => x"80", -- $09450
          37969 => x"80", -- $09451
          37970 => x"80", -- $09452
          37971 => x"80", -- $09453
          37972 => x"80", -- $09454
          37973 => x"80", -- $09455
          37974 => x"80", -- $09456
          37975 => x"80", -- $09457
          37976 => x"80", -- $09458
          37977 => x"80", -- $09459
          37978 => x"80", -- $0945a
          37979 => x"80", -- $0945b
          37980 => x"80", -- $0945c
          37981 => x"80", -- $0945d
          37982 => x"80", -- $0945e
          37983 => x"80", -- $0945f
          37984 => x"80", -- $09460
          37985 => x"80", -- $09461
          37986 => x"80", -- $09462
          37987 => x"80", -- $09463
          37988 => x"80", -- $09464
          37989 => x"80", -- $09465
          37990 => x"80", -- $09466
          37991 => x"80", -- $09467
          37992 => x"80", -- $09468
          37993 => x"80", -- $09469
          37994 => x"80", -- $0946a
          37995 => x"80", -- $0946b
          37996 => x"80", -- $0946c
          37997 => x"80", -- $0946d
          37998 => x"80", -- $0946e
          37999 => x"80", -- $0946f
          38000 => x"80", -- $09470
          38001 => x"80", -- $09471
          38002 => x"80", -- $09472
          38003 => x"80", -- $09473
          38004 => x"80", -- $09474
          38005 => x"80", -- $09475
          38006 => x"80", -- $09476
          38007 => x"80", -- $09477
          38008 => x"80", -- $09478
          38009 => x"80", -- $09479
          38010 => x"80", -- $0947a
          38011 => x"80", -- $0947b
          38012 => x"80", -- $0947c
          38013 => x"80", -- $0947d
          38014 => x"80", -- $0947e
          38015 => x"80", -- $0947f
          38016 => x"80", -- $09480
          38017 => x"80", -- $09481
          38018 => x"80", -- $09482
          38019 => x"80", -- $09483
          38020 => x"80", -- $09484
          38021 => x"80", -- $09485
          38022 => x"80", -- $09486
          38023 => x"80", -- $09487
          38024 => x"80", -- $09488
          38025 => x"80", -- $09489
          38026 => x"80", -- $0948a
          38027 => x"80", -- $0948b
          38028 => x"80", -- $0948c
          38029 => x"80", -- $0948d
          38030 => x"80", -- $0948e
          38031 => x"80", -- $0948f
          38032 => x"80", -- $09490
          38033 => x"80", -- $09491
          38034 => x"80", -- $09492
          38035 => x"80", -- $09493
          38036 => x"80", -- $09494
          38037 => x"80", -- $09495
          38038 => x"80", -- $09496
          38039 => x"80", -- $09497
          38040 => x"80", -- $09498
          38041 => x"80", -- $09499
          38042 => x"80", -- $0949a
          38043 => x"80", -- $0949b
          38044 => x"80", -- $0949c
          38045 => x"80", -- $0949d
          38046 => x"80", -- $0949e
          38047 => x"80", -- $0949f
          38048 => x"80", -- $094a0
          38049 => x"80", -- $094a1
          38050 => x"80", -- $094a2
          38051 => x"80", -- $094a3
          38052 => x"80", -- $094a4
          38053 => x"80", -- $094a5
          38054 => x"80", -- $094a6
          38055 => x"80", -- $094a7
          38056 => x"80", -- $094a8
          38057 => x"80", -- $094a9
          38058 => x"80", -- $094aa
          38059 => x"80", -- $094ab
          38060 => x"80", -- $094ac
          38061 => x"80", -- $094ad
          38062 => x"80", -- $094ae
          38063 => x"80", -- $094af
          38064 => x"80", -- $094b0
          38065 => x"80", -- $094b1
          38066 => x"80", -- $094b2
          38067 => x"80", -- $094b3
          38068 => x"80", -- $094b4
          38069 => x"80", -- $094b5
          38070 => x"80", -- $094b6
          38071 => x"80", -- $094b7
          38072 => x"80", -- $094b8
          38073 => x"80", -- $094b9
          38074 => x"80", -- $094ba
          38075 => x"80", -- $094bb
          38076 => x"80", -- $094bc
          38077 => x"80", -- $094bd
          38078 => x"80", -- $094be
          38079 => x"80", -- $094bf
          38080 => x"80", -- $094c0
          38081 => x"80", -- $094c1
          38082 => x"80", -- $094c2
          38083 => x"80", -- $094c3
          38084 => x"80", -- $094c4
          38085 => x"80", -- $094c5
          38086 => x"80", -- $094c6
          38087 => x"80", -- $094c7
          38088 => x"80", -- $094c8
          38089 => x"80", -- $094c9
          38090 => x"80", -- $094ca
          38091 => x"80", -- $094cb
          38092 => x"80", -- $094cc
          38093 => x"80", -- $094cd
          38094 => x"80", -- $094ce
          38095 => x"80", -- $094cf
          38096 => x"80", -- $094d0
          38097 => x"80", -- $094d1
          38098 => x"80", -- $094d2
          38099 => x"80", -- $094d3
          38100 => x"80", -- $094d4
          38101 => x"80", -- $094d5
          38102 => x"80", -- $094d6
          38103 => x"80", -- $094d7
          38104 => x"80", -- $094d8
          38105 => x"80", -- $094d9
          38106 => x"80", -- $094da
          38107 => x"80", -- $094db
          38108 => x"80", -- $094dc
          38109 => x"80", -- $094dd
          38110 => x"80", -- $094de
          38111 => x"80", -- $094df
          38112 => x"80", -- $094e0
          38113 => x"80", -- $094e1
          38114 => x"80", -- $094e2
          38115 => x"80", -- $094e3
          38116 => x"80", -- $094e4
          38117 => x"80", -- $094e5
          38118 => x"80", -- $094e6
          38119 => x"80", -- $094e7
          38120 => x"80", -- $094e8
          38121 => x"80", -- $094e9
          38122 => x"80", -- $094ea
          38123 => x"80", -- $094eb
          38124 => x"80", -- $094ec
          38125 => x"80", -- $094ed
          38126 => x"80", -- $094ee
          38127 => x"80", -- $094ef
          38128 => x"80", -- $094f0
          38129 => x"80", -- $094f1
          38130 => x"80", -- $094f2
          38131 => x"80", -- $094f3
          38132 => x"80", -- $094f4
          38133 => x"80", -- $094f5
          38134 => x"80", -- $094f6
          38135 => x"80", -- $094f7
          38136 => x"80", -- $094f8
          38137 => x"80", -- $094f9
          38138 => x"80", -- $094fa
          38139 => x"80", -- $094fb
          38140 => x"80", -- $094fc
          38141 => x"80", -- $094fd
          38142 => x"80", -- $094fe
          38143 => x"80", -- $094ff
          38144 => x"80", -- $09500
          38145 => x"80", -- $09501
          38146 => x"80", -- $09502
          38147 => x"80", -- $09503
          38148 => x"80", -- $09504
          38149 => x"80", -- $09505
          38150 => x"80", -- $09506
          38151 => x"80", -- $09507
          38152 => x"80", -- $09508
          38153 => x"80", -- $09509
          38154 => x"80", -- $0950a
          38155 => x"80", -- $0950b
          38156 => x"80", -- $0950c
          38157 => x"80", -- $0950d
          38158 => x"80", -- $0950e
          38159 => x"80", -- $0950f
          38160 => x"80", -- $09510
          38161 => x"80", -- $09511
          38162 => x"80", -- $09512
          38163 => x"80", -- $09513
          38164 => x"80", -- $09514
          38165 => x"80", -- $09515
          38166 => x"80", -- $09516
          38167 => x"80", -- $09517
          38168 => x"80", -- $09518
          38169 => x"80", -- $09519
          38170 => x"80", -- $0951a
          38171 => x"80", -- $0951b
          38172 => x"80", -- $0951c
          38173 => x"80", -- $0951d
          38174 => x"80", -- $0951e
          38175 => x"80", -- $0951f
          38176 => x"80", -- $09520
          38177 => x"80", -- $09521
          38178 => x"80", -- $09522
          38179 => x"80", -- $09523
          38180 => x"80", -- $09524
          38181 => x"80", -- $09525
          38182 => x"80", -- $09526
          38183 => x"80", -- $09527
          38184 => x"80", -- $09528
          38185 => x"80", -- $09529
          38186 => x"80", -- $0952a
          38187 => x"80", -- $0952b
          38188 => x"80", -- $0952c
          38189 => x"80", -- $0952d
          38190 => x"80", -- $0952e
          38191 => x"80", -- $0952f
          38192 => x"80", -- $09530
          38193 => x"80", -- $09531
          38194 => x"80", -- $09532
          38195 => x"80", -- $09533
          38196 => x"80", -- $09534
          38197 => x"80", -- $09535
          38198 => x"80", -- $09536
          38199 => x"80", -- $09537
          38200 => x"80", -- $09538
          38201 => x"80", -- $09539
          38202 => x"80", -- $0953a
          38203 => x"80", -- $0953b
          38204 => x"80", -- $0953c
          38205 => x"80", -- $0953d
          38206 => x"80", -- $0953e
          38207 => x"80", -- $0953f
          38208 => x"80", -- $09540
          38209 => x"80", -- $09541
          38210 => x"80", -- $09542
          38211 => x"80", -- $09543
          38212 => x"80", -- $09544
          38213 => x"80", -- $09545
          38214 => x"80", -- $09546
          38215 => x"80", -- $09547
          38216 => x"80", -- $09548
          38217 => x"80", -- $09549
          38218 => x"80", -- $0954a
          38219 => x"81", -- $0954b
          38220 => x"81", -- $0954c
          38221 => x"81", -- $0954d
          38222 => x"81", -- $0954e
          38223 => x"81", -- $0954f
          38224 => x"81", -- $09550
          38225 => x"81", -- $09551
          38226 => x"81", -- $09552
          38227 => x"81", -- $09553
          38228 => x"80", -- $09554
          38229 => x"80", -- $09555
          38230 => x"80", -- $09556
          38231 => x"80", -- $09557
          38232 => x"80", -- $09558
          38233 => x"80", -- $09559
          38234 => x"80", -- $0955a
          38235 => x"80", -- $0955b
          38236 => x"80", -- $0955c
          38237 => x"80", -- $0955d
          38238 => x"80", -- $0955e
          38239 => x"80", -- $0955f
          38240 => x"80", -- $09560
          38241 => x"80", -- $09561
          38242 => x"80", -- $09562
          38243 => x"80", -- $09563
          38244 => x"80", -- $09564
          38245 => x"80", -- $09565
          38246 => x"80", -- $09566
          38247 => x"80", -- $09567
          38248 => x"81", -- $09568
          38249 => x"81", -- $09569
          38250 => x"81", -- $0956a
          38251 => x"80", -- $0956b
          38252 => x"80", -- $0956c
          38253 => x"80", -- $0956d
          38254 => x"80", -- $0956e
          38255 => x"80", -- $0956f
          38256 => x"80", -- $09570
          38257 => x"80", -- $09571
          38258 => x"80", -- $09572
          38259 => x"80", -- $09573
          38260 => x"80", -- $09574
          38261 => x"80", -- $09575
          38262 => x"80", -- $09576
          38263 => x"80", -- $09577
          38264 => x"80", -- $09578
          38265 => x"80", -- $09579
          38266 => x"80", -- $0957a
          38267 => x"80", -- $0957b
          38268 => x"80", -- $0957c
          38269 => x"80", -- $0957d
          38270 => x"80", -- $0957e
          38271 => x"80", -- $0957f
          38272 => x"80", -- $09580
          38273 => x"80", -- $09581
          38274 => x"80", -- $09582
          38275 => x"80", -- $09583
          38276 => x"80", -- $09584
          38277 => x"80", -- $09585
          38278 => x"80", -- $09586
          38279 => x"80", -- $09587
          38280 => x"80", -- $09588
          38281 => x"80", -- $09589
          38282 => x"80", -- $0958a
          38283 => x"80", -- $0958b
          38284 => x"80", -- $0958c
          38285 => x"80", -- $0958d
          38286 => x"80", -- $0958e
          38287 => x"80", -- $0958f
          38288 => x"80", -- $09590
          38289 => x"80", -- $09591
          38290 => x"80", -- $09592
          38291 => x"80", -- $09593
          38292 => x"80", -- $09594
          38293 => x"80", -- $09595
          38294 => x"80", -- $09596
          38295 => x"80", -- $09597
          38296 => x"80", -- $09598
          38297 => x"80", -- $09599
          38298 => x"80", -- $0959a
          38299 => x"80", -- $0959b
          38300 => x"80", -- $0959c
          38301 => x"80", -- $0959d
          38302 => x"80", -- $0959e
          38303 => x"80", -- $0959f
          38304 => x"80", -- $095a0
          38305 => x"80", -- $095a1
          38306 => x"80", -- $095a2
          38307 => x"80", -- $095a3
          38308 => x"80", -- $095a4
          38309 => x"80", -- $095a5
          38310 => x"80", -- $095a6
          38311 => x"80", -- $095a7
          38312 => x"80", -- $095a8
          38313 => x"80", -- $095a9
          38314 => x"80", -- $095aa
          38315 => x"80", -- $095ab
          38316 => x"80", -- $095ac
          38317 => x"80", -- $095ad
          38318 => x"80", -- $095ae
          38319 => x"80", -- $095af
          38320 => x"80", -- $095b0
          38321 => x"80", -- $095b1
          38322 => x"80", -- $095b2
          38323 => x"80", -- $095b3
          38324 => x"80", -- $095b4
          38325 => x"80", -- $095b5
          38326 => x"80", -- $095b6
          38327 => x"80", -- $095b7
          38328 => x"80", -- $095b8
          38329 => x"80", -- $095b9
          38330 => x"80", -- $095ba
          38331 => x"80", -- $095bb
          38332 => x"80", -- $095bc
          38333 => x"80", -- $095bd
          38334 => x"80", -- $095be
          38335 => x"80", -- $095bf
          38336 => x"80", -- $095c0
          38337 => x"80", -- $095c1
          38338 => x"80", -- $095c2
          38339 => x"80", -- $095c3
          38340 => x"80", -- $095c4
          38341 => x"80", -- $095c5
          38342 => x"80", -- $095c6
          38343 => x"80", -- $095c7
          38344 => x"80", -- $095c8
          38345 => x"80", -- $095c9
          38346 => x"80", -- $095ca
          38347 => x"80", -- $095cb
          38348 => x"80", -- $095cc
          38349 => x"80", -- $095cd
          38350 => x"80", -- $095ce
          38351 => x"80", -- $095cf
          38352 => x"80", -- $095d0
          38353 => x"80", -- $095d1
          38354 => x"80", -- $095d2
          38355 => x"80", -- $095d3
          38356 => x"80", -- $095d4
          38357 => x"80", -- $095d5
          38358 => x"80", -- $095d6
          38359 => x"80", -- $095d7
          38360 => x"80", -- $095d8
          38361 => x"80", -- $095d9
          38362 => x"80", -- $095da
          38363 => x"80", -- $095db
          38364 => x"80", -- $095dc
          38365 => x"80", -- $095dd
          38366 => x"80", -- $095de
          38367 => x"80", -- $095df
          38368 => x"80", -- $095e0
          38369 => x"80", -- $095e1
          38370 => x"80", -- $095e2
          38371 => x"80", -- $095e3
          38372 => x"80", -- $095e4
          38373 => x"80", -- $095e5
          38374 => x"80", -- $095e6
          38375 => x"81", -- $095e7
          38376 => x"81", -- $095e8
          38377 => x"81", -- $095e9
          38378 => x"81", -- $095ea
          38379 => x"81", -- $095eb
          38380 => x"81", -- $095ec
          38381 => x"81", -- $095ed
          38382 => x"81", -- $095ee
          38383 => x"81", -- $095ef
          38384 => x"81", -- $095f0
          38385 => x"81", -- $095f1
          38386 => x"81", -- $095f2
          38387 => x"80", -- $095f3
          38388 => x"80", -- $095f4
          38389 => x"80", -- $095f5
          38390 => x"80", -- $095f6
          38391 => x"80", -- $095f7
          38392 => x"80", -- $095f8
          38393 => x"80", -- $095f9
          38394 => x"80", -- $095fa
          38395 => x"80", -- $095fb
          38396 => x"80", -- $095fc
          38397 => x"80", -- $095fd
          38398 => x"80", -- $095fe
          38399 => x"80", -- $095ff
          38400 => x"80", -- $09600
          38401 => x"80", -- $09601
          38402 => x"81", -- $09602
          38403 => x"81", -- $09603
          38404 => x"81", -- $09604
          38405 => x"81", -- $09605
          38406 => x"81", -- $09606
          38407 => x"81", -- $09607
          38408 => x"81", -- $09608
          38409 => x"81", -- $09609
          38410 => x"81", -- $0960a
          38411 => x"81", -- $0960b
          38412 => x"81", -- $0960c
          38413 => x"81", -- $0960d
          38414 => x"81", -- $0960e
          38415 => x"81", -- $0960f
          38416 => x"81", -- $09610
          38417 => x"80", -- $09611
          38418 => x"80", -- $09612
          38419 => x"80", -- $09613
          38420 => x"80", -- $09614
          38421 => x"80", -- $09615
          38422 => x"80", -- $09616
          38423 => x"80", -- $09617
          38424 => x"80", -- $09618
          38425 => x"80", -- $09619
          38426 => x"80", -- $0961a
          38427 => x"80", -- $0961b
          38428 => x"80", -- $0961c
          38429 => x"80", -- $0961d
          38430 => x"80", -- $0961e
          38431 => x"80", -- $0961f
          38432 => x"80", -- $09620
          38433 => x"80", -- $09621
          38434 => x"80", -- $09622
          38435 => x"80", -- $09623
          38436 => x"80", -- $09624
          38437 => x"80", -- $09625
          38438 => x"80", -- $09626
          38439 => x"80", -- $09627
          38440 => x"80", -- $09628
          38441 => x"80", -- $09629
          38442 => x"80", -- $0962a
          38443 => x"80", -- $0962b
          38444 => x"80", -- $0962c
          38445 => x"80", -- $0962d
          38446 => x"80", -- $0962e
          38447 => x"80", -- $0962f
          38448 => x"80", -- $09630
          38449 => x"80", -- $09631
          38450 => x"80", -- $09632
          38451 => x"80", -- $09633
          38452 => x"80", -- $09634
          38453 => x"80", -- $09635
          38454 => x"80", -- $09636
          38455 => x"80", -- $09637
          38456 => x"80", -- $09638
          38457 => x"80", -- $09639
          38458 => x"80", -- $0963a
          38459 => x"80", -- $0963b
          38460 => x"80", -- $0963c
          38461 => x"80", -- $0963d
          38462 => x"80", -- $0963e
          38463 => x"80", -- $0963f
          38464 => x"80", -- $09640
          38465 => x"80", -- $09641
          38466 => x"80", -- $09642
          38467 => x"80", -- $09643
          38468 => x"80", -- $09644
          38469 => x"80", -- $09645
          38470 => x"80", -- $09646
          38471 => x"80", -- $09647
          38472 => x"80", -- $09648
          38473 => x"80", -- $09649
          38474 => x"80", -- $0964a
          38475 => x"80", -- $0964b
          38476 => x"80", -- $0964c
          38477 => x"80", -- $0964d
          38478 => x"80", -- $0964e
          38479 => x"80", -- $0964f
          38480 => x"80", -- $09650
          38481 => x"80", -- $09651
          38482 => x"80", -- $09652
          38483 => x"80", -- $09653
          38484 => x"80", -- $09654
          38485 => x"80", -- $09655
          38486 => x"80", -- $09656
          38487 => x"80", -- $09657
          38488 => x"80", -- $09658
          38489 => x"80", -- $09659
          38490 => x"80", -- $0965a
          38491 => x"80", -- $0965b
          38492 => x"80", -- $0965c
          38493 => x"80", -- $0965d
          38494 => x"80", -- $0965e
          38495 => x"80", -- $0965f
          38496 => x"80", -- $09660
          38497 => x"80", -- $09661
          38498 => x"80", -- $09662
          38499 => x"80", -- $09663
          38500 => x"80", -- $09664
          38501 => x"80", -- $09665
          38502 => x"80", -- $09666
          38503 => x"80", -- $09667
          38504 => x"80", -- $09668
          38505 => x"80", -- $09669
          38506 => x"80", -- $0966a
          38507 => x"80", -- $0966b
          38508 => x"80", -- $0966c
          38509 => x"80", -- $0966d
          38510 => x"80", -- $0966e
          38511 => x"80", -- $0966f
          38512 => x"80", -- $09670
          38513 => x"80", -- $09671
          38514 => x"80", -- $09672
          38515 => x"80", -- $09673
          38516 => x"80", -- $09674
          38517 => x"80", -- $09675
          38518 => x"7f", -- $09676
          38519 => x"7f", -- $09677
          38520 => x"7f", -- $09678
          38521 => x"80", -- $09679
          38522 => x"7f", -- $0967a
          38523 => x"7f", -- $0967b
          38524 => x"7f", -- $0967c
          38525 => x"7f", -- $0967d
          38526 => x"7f", -- $0967e
          38527 => x"7f", -- $0967f
          38528 => x"80", -- $09680
          38529 => x"80", -- $09681
          38530 => x"80", -- $09682
          38531 => x"80", -- $09683
          38532 => x"80", -- $09684
          38533 => x"80", -- $09685
          38534 => x"80", -- $09686
          38535 => x"80", -- $09687
          38536 => x"80", -- $09688
          38537 => x"80", -- $09689
          38538 => x"80", -- $0968a
          38539 => x"80", -- $0968b
          38540 => x"80", -- $0968c
          38541 => x"80", -- $0968d
          38542 => x"80", -- $0968e
          38543 => x"80", -- $0968f
          38544 => x"80", -- $09690
          38545 => x"80", -- $09691
          38546 => x"80", -- $09692
          38547 => x"80", -- $09693
          38548 => x"80", -- $09694
          38549 => x"80", -- $09695
          38550 => x"7f", -- $09696
          38551 => x"7f", -- $09697
          38552 => x"7f", -- $09698
          38553 => x"7f", -- $09699
          38554 => x"7f", -- $0969a
          38555 => x"7f", -- $0969b
          38556 => x"7f", -- $0969c
          38557 => x"7f", -- $0969d
          38558 => x"80", -- $0969e
          38559 => x"80", -- $0969f
          38560 => x"80", -- $096a0
          38561 => x"80", -- $096a1
          38562 => x"80", -- $096a2
          38563 => x"80", -- $096a3
          38564 => x"80", -- $096a4
          38565 => x"80", -- $096a5
          38566 => x"80", -- $096a6
          38567 => x"80", -- $096a7
          38568 => x"80", -- $096a8
          38569 => x"80", -- $096a9
          38570 => x"80", -- $096aa
          38571 => x"80", -- $096ab
          38572 => x"80", -- $096ac
          38573 => x"80", -- $096ad
          38574 => x"80", -- $096ae
          38575 => x"80", -- $096af
          38576 => x"80", -- $096b0
          38577 => x"80", -- $096b1
          38578 => x"80", -- $096b2
          38579 => x"80", -- $096b3
          38580 => x"80", -- $096b4
          38581 => x"80", -- $096b5
          38582 => x"80", -- $096b6
          38583 => x"80", -- $096b7
          38584 => x"80", -- $096b8
          38585 => x"80", -- $096b9
          38586 => x"80", -- $096ba
          38587 => x"80", -- $096bb
          38588 => x"80", -- $096bc
          38589 => x"80", -- $096bd
          38590 => x"80", -- $096be
          38591 => x"80", -- $096bf
          38592 => x"80", -- $096c0
          38593 => x"80", -- $096c1
          38594 => x"80", -- $096c2
          38595 => x"80", -- $096c3
          38596 => x"80", -- $096c4
          38597 => x"80", -- $096c5
          38598 => x"80", -- $096c6
          38599 => x"80", -- $096c7
          38600 => x"80", -- $096c8
          38601 => x"80", -- $096c9
          38602 => x"80", -- $096ca
          38603 => x"80", -- $096cb
          38604 => x"80", -- $096cc
          38605 => x"80", -- $096cd
          38606 => x"80", -- $096ce
          38607 => x"80", -- $096cf
          38608 => x"80", -- $096d0
          38609 => x"80", -- $096d1
          38610 => x"80", -- $096d2
          38611 => x"80", -- $096d3
          38612 => x"80", -- $096d4
          38613 => x"80", -- $096d5
          38614 => x"80", -- $096d6
          38615 => x"80", -- $096d7
          38616 => x"80", -- $096d8
          38617 => x"80", -- $096d9
          38618 => x"80", -- $096da
          38619 => x"80", -- $096db
          38620 => x"80", -- $096dc
          38621 => x"80", -- $096dd
          38622 => x"80", -- $096de
          38623 => x"80", -- $096df
          38624 => x"80", -- $096e0
          38625 => x"80", -- $096e1
          38626 => x"80", -- $096e2
          38627 => x"80", -- $096e3
          38628 => x"80", -- $096e4
          38629 => x"80", -- $096e5
          38630 => x"80", -- $096e6
          38631 => x"80", -- $096e7
          38632 => x"80", -- $096e8
          38633 => x"80", -- $096e9
          38634 => x"80", -- $096ea
          38635 => x"80", -- $096eb
          38636 => x"80", -- $096ec
          38637 => x"80", -- $096ed
          38638 => x"80", -- $096ee
          38639 => x"80", -- $096ef
          38640 => x"80", -- $096f0
          38641 => x"80", -- $096f1
          38642 => x"80", -- $096f2
          38643 => x"80", -- $096f3
          38644 => x"80", -- $096f4
          38645 => x"80", -- $096f5
          38646 => x"80", -- $096f6
          38647 => x"80", -- $096f7
          38648 => x"80", -- $096f8
          38649 => x"80", -- $096f9
          38650 => x"80", -- $096fa
          38651 => x"80", -- $096fb
          38652 => x"80", -- $096fc
          38653 => x"80", -- $096fd
          38654 => x"80", -- $096fe
          38655 => x"80", -- $096ff
          38656 => x"80", -- $09700
          38657 => x"80", -- $09701
          38658 => x"80", -- $09702
          38659 => x"80", -- $09703
          38660 => x"80", -- $09704
          38661 => x"80", -- $09705
          38662 => x"80", -- $09706
          38663 => x"80", -- $09707
          38664 => x"80", -- $09708
          38665 => x"80", -- $09709
          38666 => x"80", -- $0970a
          38667 => x"80", -- $0970b
          38668 => x"80", -- $0970c
          38669 => x"80", -- $0970d
          38670 => x"80", -- $0970e
          38671 => x"80", -- $0970f
          38672 => x"80", -- $09710
          38673 => x"80", -- $09711
          38674 => x"80", -- $09712
          38675 => x"80", -- $09713
          38676 => x"80", -- $09714
          38677 => x"80", -- $09715
          38678 => x"80", -- $09716
          38679 => x"80", -- $09717
          38680 => x"80", -- $09718
          38681 => x"80", -- $09719
          38682 => x"80", -- $0971a
          38683 => x"80", -- $0971b
          38684 => x"80", -- $0971c
          38685 => x"80", -- $0971d
          38686 => x"80", -- $0971e
          38687 => x"80", -- $0971f
          38688 => x"80", -- $09720
          38689 => x"80", -- $09721
          38690 => x"80", -- $09722
          38691 => x"80", -- $09723
          38692 => x"80", -- $09724
          38693 => x"80", -- $09725
          38694 => x"80", -- $09726
          38695 => x"80", -- $09727
          38696 => x"80", -- $09728
          38697 => x"80", -- $09729
          38698 => x"80", -- $0972a
          38699 => x"80", -- $0972b
          38700 => x"80", -- $0972c
          38701 => x"80", -- $0972d
          38702 => x"80", -- $0972e
          38703 => x"80", -- $0972f
          38704 => x"80", -- $09730
          38705 => x"80", -- $09731
          38706 => x"80", -- $09732
          38707 => x"80", -- $09733
          38708 => x"80", -- $09734
          38709 => x"80", -- $09735
          38710 => x"80", -- $09736
          38711 => x"80", -- $09737
          38712 => x"80", -- $09738
          38713 => x"80", -- $09739
          38714 => x"80", -- $0973a
          38715 => x"80", -- $0973b
          38716 => x"80", -- $0973c
          38717 => x"80", -- $0973d
          38718 => x"80", -- $0973e
          38719 => x"80", -- $0973f
          38720 => x"80", -- $09740
          38721 => x"80", -- $09741
          38722 => x"80", -- $09742
          38723 => x"80", -- $09743
          38724 => x"80", -- $09744
          38725 => x"80", -- $09745
          38726 => x"80", -- $09746
          38727 => x"80", -- $09747
          38728 => x"80", -- $09748
          38729 => x"80", -- $09749
          38730 => x"80", -- $0974a
          38731 => x"80", -- $0974b
          38732 => x"80", -- $0974c
          38733 => x"80", -- $0974d
          38734 => x"80", -- $0974e
          38735 => x"80", -- $0974f
          38736 => x"80", -- $09750
          38737 => x"80", -- $09751
          38738 => x"80", -- $09752
          38739 => x"80", -- $09753
          38740 => x"80", -- $09754
          38741 => x"80", -- $09755
          38742 => x"80", -- $09756
          38743 => x"80", -- $09757
          38744 => x"80", -- $09758
          38745 => x"80", -- $09759
          38746 => x"80", -- $0975a
          38747 => x"80", -- $0975b
          38748 => x"80", -- $0975c
          38749 => x"80", -- $0975d
          38750 => x"80", -- $0975e
          38751 => x"80", -- $0975f
          38752 => x"80", -- $09760
          38753 => x"80", -- $09761
          38754 => x"80", -- $09762
          38755 => x"80", -- $09763
          38756 => x"80", -- $09764
          38757 => x"80", -- $09765
          38758 => x"80", -- $09766
          38759 => x"80", -- $09767
          38760 => x"80", -- $09768
          38761 => x"80", -- $09769
          38762 => x"80", -- $0976a
          38763 => x"80", -- $0976b
          38764 => x"80", -- $0976c
          38765 => x"80", -- $0976d
          38766 => x"80", -- $0976e
          38767 => x"80", -- $0976f
          38768 => x"80", -- $09770
          38769 => x"80", -- $09771
          38770 => x"80", -- $09772
          38771 => x"80", -- $09773
          38772 => x"80", -- $09774
          38773 => x"80", -- $09775
          38774 => x"80", -- $09776
          38775 => x"80", -- $09777
          38776 => x"80", -- $09778
          38777 => x"80", -- $09779
          38778 => x"80", -- $0977a
          38779 => x"80", -- $0977b
          38780 => x"80", -- $0977c
          38781 => x"80", -- $0977d
          38782 => x"80", -- $0977e
          38783 => x"80", -- $0977f
          38784 => x"80", -- $09780
          38785 => x"80", -- $09781
          38786 => x"80", -- $09782
          38787 => x"80", -- $09783
          38788 => x"80", -- $09784
          38789 => x"80", -- $09785
          38790 => x"80", -- $09786
          38791 => x"80", -- $09787
          38792 => x"80", -- $09788
          38793 => x"80", -- $09789
          38794 => x"80", -- $0978a
          38795 => x"80", -- $0978b
          38796 => x"80", -- $0978c
          38797 => x"80", -- $0978d
          38798 => x"80", -- $0978e
          38799 => x"80", -- $0978f
          38800 => x"80", -- $09790
          38801 => x"80", -- $09791
          38802 => x"80", -- $09792
          38803 => x"80", -- $09793
          38804 => x"80", -- $09794
          38805 => x"80", -- $09795
          38806 => x"80", -- $09796
          38807 => x"80", -- $09797
          38808 => x"80", -- $09798
          38809 => x"80", -- $09799
          38810 => x"80", -- $0979a
          38811 => x"80", -- $0979b
          38812 => x"80", -- $0979c
          38813 => x"80", -- $0979d
          38814 => x"80", -- $0979e
          38815 => x"80", -- $0979f
          38816 => x"80", -- $097a0
          38817 => x"80", -- $097a1
          38818 => x"80", -- $097a2
          38819 => x"80", -- $097a3
          38820 => x"80", -- $097a4
          38821 => x"80", -- $097a5
          38822 => x"80", -- $097a6
          38823 => x"80", -- $097a7
          38824 => x"80", -- $097a8
          38825 => x"80", -- $097a9
          38826 => x"80", -- $097aa
          38827 => x"80", -- $097ab
          38828 => x"80", -- $097ac
          38829 => x"80", -- $097ad
          38830 => x"80", -- $097ae
          38831 => x"80", -- $097af
          38832 => x"80", -- $097b0
          38833 => x"80", -- $097b1
          38834 => x"80", -- $097b2
          38835 => x"80", -- $097b3
          38836 => x"80", -- $097b4
          38837 => x"80", -- $097b5
          38838 => x"80", -- $097b6
          38839 => x"80", -- $097b7
          38840 => x"80", -- $097b8
          38841 => x"80", -- $097b9
          38842 => x"80", -- $097ba
          38843 => x"80", -- $097bb
          38844 => x"80", -- $097bc
          38845 => x"80", -- $097bd
          38846 => x"80", -- $097be
          38847 => x"80", -- $097bf
          38848 => x"80", -- $097c0
          38849 => x"80", -- $097c1
          38850 => x"80", -- $097c2
          38851 => x"80", -- $097c3
          38852 => x"80", -- $097c4
          38853 => x"80", -- $097c5
          38854 => x"80", -- $097c6
          38855 => x"80", -- $097c7
          38856 => x"80", -- $097c8
          38857 => x"80", -- $097c9
          38858 => x"80", -- $097ca
          38859 => x"80", -- $097cb
          38860 => x"80", -- $097cc
          38861 => x"81", -- $097cd
          38862 => x"80", -- $097ce
          38863 => x"80", -- $097cf
          38864 => x"80", -- $097d0
          38865 => x"81", -- $097d1
          38866 => x"80", -- $097d2
          38867 => x"80", -- $097d3
          38868 => x"80", -- $097d4
          38869 => x"80", -- $097d5
          38870 => x"80", -- $097d6
          38871 => x"80", -- $097d7
          38872 => x"80", -- $097d8
          38873 => x"80", -- $097d9
          38874 => x"80", -- $097da
          38875 => x"80", -- $097db
          38876 => x"80", -- $097dc
          38877 => x"80", -- $097dd
          38878 => x"80", -- $097de
          38879 => x"80", -- $097df
          38880 => x"80", -- $097e0
          38881 => x"80", -- $097e1
          38882 => x"80", -- $097e2
          38883 => x"80", -- $097e3
          38884 => x"80", -- $097e4
          38885 => x"80", -- $097e5
          38886 => x"80", -- $097e6
          38887 => x"80", -- $097e7
          38888 => x"80", -- $097e8
          38889 => x"80", -- $097e9
          38890 => x"80", -- $097ea
          38891 => x"80", -- $097eb
          38892 => x"80", -- $097ec
          38893 => x"80", -- $097ed
          38894 => x"80", -- $097ee
          38895 => x"80", -- $097ef
          38896 => x"80", -- $097f0
          38897 => x"80", -- $097f1
          38898 => x"80", -- $097f2
          38899 => x"80", -- $097f3
          38900 => x"80", -- $097f4
          38901 => x"80", -- $097f5
          38902 => x"80", -- $097f6
          38903 => x"80", -- $097f7
          38904 => x"80", -- $097f8
          38905 => x"80", -- $097f9
          38906 => x"80", -- $097fa
          38907 => x"80", -- $097fb
          38908 => x"80", -- $097fc
          38909 => x"80", -- $097fd
          38910 => x"80", -- $097fe
          38911 => x"80", -- $097ff
          38912 => x"80", -- $09800
          38913 => x"80", -- $09801
          38914 => x"80", -- $09802
          38915 => x"80", -- $09803
          38916 => x"80", -- $09804
          38917 => x"80", -- $09805
          38918 => x"80", -- $09806
          38919 => x"80", -- $09807
          38920 => x"80", -- $09808
          38921 => x"80", -- $09809
          38922 => x"80", -- $0980a
          38923 => x"80", -- $0980b
          38924 => x"80", -- $0980c
          38925 => x"80", -- $0980d
          38926 => x"80", -- $0980e
          38927 => x"80", -- $0980f
          38928 => x"80", -- $09810
          38929 => x"80", -- $09811
          38930 => x"80", -- $09812
          38931 => x"80", -- $09813
          38932 => x"80", -- $09814
          38933 => x"80", -- $09815
          38934 => x"80", -- $09816
          38935 => x"80", -- $09817
          38936 => x"80", -- $09818
          38937 => x"80", -- $09819
          38938 => x"80", -- $0981a
          38939 => x"80", -- $0981b
          38940 => x"80", -- $0981c
          38941 => x"80", -- $0981d
          38942 => x"80", -- $0981e
          38943 => x"80", -- $0981f
          38944 => x"80", -- $09820
          38945 => x"80", -- $09821
          38946 => x"80", -- $09822
          38947 => x"80", -- $09823
          38948 => x"80", -- $09824
          38949 => x"80", -- $09825
          38950 => x"80", -- $09826
          38951 => x"80", -- $09827
          38952 => x"80", -- $09828
          38953 => x"80", -- $09829
          38954 => x"80", -- $0982a
          38955 => x"80", -- $0982b
          38956 => x"80", -- $0982c
          38957 => x"80", -- $0982d
          38958 => x"80", -- $0982e
          38959 => x"80", -- $0982f
          38960 => x"80", -- $09830
          38961 => x"80", -- $09831
          38962 => x"80", -- $09832
          38963 => x"80", -- $09833
          38964 => x"80", -- $09834
          38965 => x"80", -- $09835
          38966 => x"80", -- $09836
          38967 => x"80", -- $09837
          38968 => x"80", -- $09838
          38969 => x"80", -- $09839
          38970 => x"80", -- $0983a
          38971 => x"80", -- $0983b
          38972 => x"80", -- $0983c
          38973 => x"80", -- $0983d
          38974 => x"80", -- $0983e
          38975 => x"80", -- $0983f
          38976 => x"80", -- $09840
          38977 => x"80", -- $09841
          38978 => x"80", -- $09842
          38979 => x"80", -- $09843
          38980 => x"80", -- $09844
          38981 => x"80", -- $09845
          38982 => x"80", -- $09846
          38983 => x"80", -- $09847
          38984 => x"80", -- $09848
          38985 => x"80", -- $09849
          38986 => x"80", -- $0984a
          38987 => x"80", -- $0984b
          38988 => x"80", -- $0984c
          38989 => x"80", -- $0984d
          38990 => x"81", -- $0984e
          38991 => x"81", -- $0984f
          38992 => x"81", -- $09850
          38993 => x"81", -- $09851
          38994 => x"81", -- $09852
          38995 => x"81", -- $09853
          38996 => x"81", -- $09854
          38997 => x"81", -- $09855
          38998 => x"81", -- $09856
          38999 => x"80", -- $09857
          39000 => x"80", -- $09858
          39001 => x"80", -- $09859
          39002 => x"80", -- $0985a
          39003 => x"80", -- $0985b
          39004 => x"80", -- $0985c
          39005 => x"80", -- $0985d
          39006 => x"80", -- $0985e
          39007 => x"80", -- $0985f
          39008 => x"80", -- $09860
          39009 => x"80", -- $09861
          39010 => x"80", -- $09862
          39011 => x"80", -- $09863
          39012 => x"80", -- $09864
          39013 => x"80", -- $09865
          39014 => x"80", -- $09866
          39015 => x"80", -- $09867
          39016 => x"80", -- $09868
          39017 => x"80", -- $09869
          39018 => x"81", -- $0986a
          39019 => x"81", -- $0986b
          39020 => x"81", -- $0986c
          39021 => x"81", -- $0986d
          39022 => x"81", -- $0986e
          39023 => x"81", -- $0986f
          39024 => x"81", -- $09870
          39025 => x"81", -- $09871
          39026 => x"81", -- $09872
          39027 => x"81", -- $09873
          39028 => x"81", -- $09874
          39029 => x"81", -- $09875
          39030 => x"81", -- $09876
          39031 => x"81", -- $09877
          39032 => x"81", -- $09878
          39033 => x"81", -- $09879
          39034 => x"81", -- $0987a
          39035 => x"81", -- $0987b
          39036 => x"80", -- $0987c
          39037 => x"80", -- $0987d
          39038 => x"80", -- $0987e
          39039 => x"80", -- $0987f
          39040 => x"80", -- $09880
          39041 => x"80", -- $09881
          39042 => x"80", -- $09882
          39043 => x"80", -- $09883
          39044 => x"80", -- $09884
          39045 => x"80", -- $09885
          39046 => x"80", -- $09886
          39047 => x"80", -- $09887
          39048 => x"80", -- $09888
          39049 => x"81", -- $09889
          39050 => x"81", -- $0988a
          39051 => x"81", -- $0988b
          39052 => x"81", -- $0988c
          39053 => x"81", -- $0988d
          39054 => x"81", -- $0988e
          39055 => x"81", -- $0988f
          39056 => x"81", -- $09890
          39057 => x"81", -- $09891
          39058 => x"81", -- $09892
          39059 => x"81", -- $09893
          39060 => x"81", -- $09894
          39061 => x"81", -- $09895
          39062 => x"81", -- $09896
          39063 => x"81", -- $09897
          39064 => x"81", -- $09898
          39065 => x"81", -- $09899
          39066 => x"81", -- $0989a
          39067 => x"81", -- $0989b
          39068 => x"81", -- $0989c
          39069 => x"81", -- $0989d
          39070 => x"80", -- $0989e
          39071 => x"80", -- $0989f
          39072 => x"80", -- $098a0
          39073 => x"80", -- $098a1
          39074 => x"80", -- $098a2
          39075 => x"80", -- $098a3
          39076 => x"80", -- $098a4
          39077 => x"80", -- $098a5
          39078 => x"80", -- $098a6
          39079 => x"80", -- $098a7
          39080 => x"80", -- $098a8
          39081 => x"80", -- $098a9
          39082 => x"80", -- $098aa
          39083 => x"81", -- $098ab
          39084 => x"81", -- $098ac
          39085 => x"81", -- $098ad
          39086 => x"81", -- $098ae
          39087 => x"81", -- $098af
          39088 => x"81", -- $098b0
          39089 => x"81", -- $098b1
          39090 => x"81", -- $098b2
          39091 => x"81", -- $098b3
          39092 => x"81", -- $098b4
          39093 => x"81", -- $098b5
          39094 => x"81", -- $098b6
          39095 => x"81", -- $098b7
          39096 => x"81", -- $098b8
          39097 => x"81", -- $098b9
          39098 => x"80", -- $098ba
          39099 => x"80", -- $098bb
          39100 => x"80", -- $098bc
          39101 => x"80", -- $098bd
          39102 => x"80", -- $098be
          39103 => x"80", -- $098bf
          39104 => x"80", -- $098c0
          39105 => x"80", -- $098c1
          39106 => x"80", -- $098c2
          39107 => x"80", -- $098c3
          39108 => x"80", -- $098c4
          39109 => x"80", -- $098c5
          39110 => x"80", -- $098c6
          39111 => x"80", -- $098c7
          39112 => x"80", -- $098c8
          39113 => x"80", -- $098c9
          39114 => x"80", -- $098ca
          39115 => x"80", -- $098cb
          39116 => x"80", -- $098cc
          39117 => x"80", -- $098cd
          39118 => x"80", -- $098ce
          39119 => x"81", -- $098cf
          39120 => x"81", -- $098d0
          39121 => x"81", -- $098d1
          39122 => x"80", -- $098d2
          39123 => x"80", -- $098d3
          39124 => x"80", -- $098d4
          39125 => x"80", -- $098d5
          39126 => x"80", -- $098d6
          39127 => x"80", -- $098d7
          39128 => x"80", -- $098d8
          39129 => x"80", -- $098d9
          39130 => x"80", -- $098da
          39131 => x"80", -- $098db
          39132 => x"80", -- $098dc
          39133 => x"80", -- $098dd
          39134 => x"80", -- $098de
          39135 => x"80", -- $098df
          39136 => x"80", -- $098e0
          39137 => x"80", -- $098e1
          39138 => x"80", -- $098e2
          39139 => x"80", -- $098e3
          39140 => x"80", -- $098e4
          39141 => x"80", -- $098e5
          39142 => x"80", -- $098e6
          39143 => x"80", -- $098e7
          39144 => x"80", -- $098e8
          39145 => x"80", -- $098e9
          39146 => x"80", -- $098ea
          39147 => x"80", -- $098eb
          39148 => x"80", -- $098ec
          39149 => x"80", -- $098ed
          39150 => x"80", -- $098ee
          39151 => x"80", -- $098ef
          39152 => x"80", -- $098f0
          39153 => x"80", -- $098f1
          39154 => x"80", -- $098f2
          39155 => x"80", -- $098f3
          39156 => x"80", -- $098f4
          39157 => x"80", -- $098f5
          39158 => x"80", -- $098f6
          39159 => x"80", -- $098f7
          39160 => x"80", -- $098f8
          39161 => x"80", -- $098f9
          39162 => x"80", -- $098fa
          39163 => x"80", -- $098fb
          39164 => x"80", -- $098fc
          39165 => x"80", -- $098fd
          39166 => x"80", -- $098fe
          39167 => x"80", -- $098ff
          39168 => x"80", -- $09900
          39169 => x"80", -- $09901
          39170 => x"80", -- $09902
          39171 => x"80", -- $09903
          39172 => x"80", -- $09904
          39173 => x"80", -- $09905
          39174 => x"80", -- $09906
          39175 => x"80", -- $09907
          39176 => x"80", -- $09908
          39177 => x"80", -- $09909
          39178 => x"80", -- $0990a
          39179 => x"80", -- $0990b
          39180 => x"80", -- $0990c
          39181 => x"80", -- $0990d
          39182 => x"80", -- $0990e
          39183 => x"80", -- $0990f
          39184 => x"80", -- $09910
          39185 => x"80", -- $09911
          39186 => x"80", -- $09912
          39187 => x"80", -- $09913
          39188 => x"80", -- $09914
          39189 => x"80", -- $09915
          39190 => x"80", -- $09916
          39191 => x"80", -- $09917
          39192 => x"80", -- $09918
          39193 => x"80", -- $09919
          39194 => x"80", -- $0991a
          39195 => x"80", -- $0991b
          39196 => x"80", -- $0991c
          39197 => x"80", -- $0991d
          39198 => x"80", -- $0991e
          39199 => x"80", -- $0991f
          39200 => x"80", -- $09920
          39201 => x"80", -- $09921
          39202 => x"80", -- $09922
          39203 => x"80", -- $09923
          39204 => x"80", -- $09924
          39205 => x"80", -- $09925
          39206 => x"80", -- $09926
          39207 => x"80", -- $09927
          39208 => x"80", -- $09928
          39209 => x"80", -- $09929
          39210 => x"80", -- $0992a
          39211 => x"80", -- $0992b
          39212 => x"80", -- $0992c
          39213 => x"80", -- $0992d
          39214 => x"80", -- $0992e
          39215 => x"80", -- $0992f
          39216 => x"80", -- $09930
          39217 => x"80", -- $09931
          39218 => x"80", -- $09932
          39219 => x"80", -- $09933
          39220 => x"80", -- $09934
          39221 => x"80", -- $09935
          39222 => x"80", -- $09936
          39223 => x"80", -- $09937
          39224 => x"80", -- $09938
          39225 => x"80", -- $09939
          39226 => x"80", -- $0993a
          39227 => x"80", -- $0993b
          39228 => x"80", -- $0993c
          39229 => x"80", -- $0993d
          39230 => x"80", -- $0993e
          39231 => x"80", -- $0993f
          39232 => x"80", -- $09940
          39233 => x"7f", -- $09941
          39234 => x"7f", -- $09942
          39235 => x"80", -- $09943
          39236 => x"80", -- $09944
          39237 => x"80", -- $09945
          39238 => x"80", -- $09946
          39239 => x"80", -- $09947
          39240 => x"80", -- $09948
          39241 => x"80", -- $09949
          39242 => x"80", -- $0994a
          39243 => x"80", -- $0994b
          39244 => x"80", -- $0994c
          39245 => x"80", -- $0994d
          39246 => x"80", -- $0994e
          39247 => x"80", -- $0994f
          39248 => x"80", -- $09950
          39249 => x"80", -- $09951
          39250 => x"80", -- $09952
          39251 => x"80", -- $09953
          39252 => x"80", -- $09954
          39253 => x"80", -- $09955
          39254 => x"80", -- $09956
          39255 => x"80", -- $09957
          39256 => x"80", -- $09958
          39257 => x"80", -- $09959
          39258 => x"80", -- $0995a
          39259 => x"80", -- $0995b
          39260 => x"80", -- $0995c
          39261 => x"80", -- $0995d
          39262 => x"80", -- $0995e
          39263 => x"80", -- $0995f
          39264 => x"80", -- $09960
          39265 => x"80", -- $09961
          39266 => x"80", -- $09962
          39267 => x"80", -- $09963
          39268 => x"80", -- $09964
          39269 => x"7f", -- $09965
          39270 => x"80", -- $09966
          39271 => x"80", -- $09967
          39272 => x"80", -- $09968
          39273 => x"80", -- $09969
          39274 => x"80", -- $0996a
          39275 => x"80", -- $0996b
          39276 => x"80", -- $0996c
          39277 => x"80", -- $0996d
          39278 => x"80", -- $0996e
          39279 => x"80", -- $0996f
          39280 => x"80", -- $09970
          39281 => x"80", -- $09971
          39282 => x"80", -- $09972
          39283 => x"80", -- $09973
          39284 => x"80", -- $09974
          39285 => x"80", -- $09975
          39286 => x"80", -- $09976
          39287 => x"80", -- $09977
          39288 => x"80", -- $09978
          39289 => x"80", -- $09979
          39290 => x"80", -- $0997a
          39291 => x"80", -- $0997b
          39292 => x"80", -- $0997c
          39293 => x"80", -- $0997d
          39294 => x"7f", -- $0997e
          39295 => x"7f", -- $0997f
          39296 => x"7f", -- $09980
          39297 => x"7f", -- $09981
          39298 => x"7f", -- $09982
          39299 => x"7f", -- $09983
          39300 => x"7f", -- $09984
          39301 => x"7f", -- $09985
          39302 => x"80", -- $09986
          39303 => x"80", -- $09987
          39304 => x"80", -- $09988
          39305 => x"80", -- $09989
          39306 => x"80", -- $0998a
          39307 => x"80", -- $0998b
          39308 => x"80", -- $0998c
          39309 => x"80", -- $0998d
          39310 => x"80", -- $0998e
          39311 => x"80", -- $0998f
          39312 => x"80", -- $09990
          39313 => x"80", -- $09991
          39314 => x"80", -- $09992
          39315 => x"80", -- $09993
          39316 => x"80", -- $09994
          39317 => x"80", -- $09995
          39318 => x"80", -- $09996
          39319 => x"80", -- $09997
          39320 => x"80", -- $09998
          39321 => x"80", -- $09999
          39322 => x"80", -- $0999a
          39323 => x"80", -- $0999b
          39324 => x"80", -- $0999c
          39325 => x"80", -- $0999d
          39326 => x"80", -- $0999e
          39327 => x"80", -- $0999f
          39328 => x"80", -- $099a0
          39329 => x"80", -- $099a1
          39330 => x"80", -- $099a2
          39331 => x"80", -- $099a3
          39332 => x"80", -- $099a4
          39333 => x"80", -- $099a5
          39334 => x"80", -- $099a6
          39335 => x"80", -- $099a7
          39336 => x"80", -- $099a8
          39337 => x"80", -- $099a9
          39338 => x"80", -- $099aa
          39339 => x"80", -- $099ab
          39340 => x"80", -- $099ac
          39341 => x"80", -- $099ad
          39342 => x"80", -- $099ae
          39343 => x"80", -- $099af
          39344 => x"80", -- $099b0
          39345 => x"80", -- $099b1
          39346 => x"80", -- $099b2
          39347 => x"80", -- $099b3
          39348 => x"80", -- $099b4
          39349 => x"80", -- $099b5
          39350 => x"80", -- $099b6
          39351 => x"80", -- $099b7
          39352 => x"80", -- $099b8
          39353 => x"80", -- $099b9
          39354 => x"80", -- $099ba
          39355 => x"80", -- $099bb
          39356 => x"80", -- $099bc
          39357 => x"80", -- $099bd
          39358 => x"80", -- $099be
          39359 => x"80", -- $099bf
          39360 => x"80", -- $099c0
          39361 => x"80", -- $099c1
          39362 => x"7f", -- $099c2
          39363 => x"7f", -- $099c3
          39364 => x"7f", -- $099c4
          39365 => x"80", -- $099c5
          39366 => x"80", -- $099c6
          39367 => x"80", -- $099c7
          39368 => x"80", -- $099c8
          39369 => x"80", -- $099c9
          39370 => x"80", -- $099ca
          39371 => x"80", -- $099cb
          39372 => x"80", -- $099cc
          39373 => x"80", -- $099cd
          39374 => x"80", -- $099ce
          39375 => x"80", -- $099cf
          39376 => x"80", -- $099d0
          39377 => x"80", -- $099d1
          39378 => x"80", -- $099d2
          39379 => x"80", -- $099d3
          39380 => x"80", -- $099d4
          39381 => x"80", -- $099d5
          39382 => x"80", -- $099d6
          39383 => x"80", -- $099d7
          39384 => x"80", -- $099d8
          39385 => x"80", -- $099d9
          39386 => x"80", -- $099da
          39387 => x"7f", -- $099db
          39388 => x"7f", -- $099dc
          39389 => x"7f", -- $099dd
          39390 => x"7f", -- $099de
          39391 => x"7f", -- $099df
          39392 => x"7f", -- $099e0
          39393 => x"7f", -- $099e1
          39394 => x"7f", -- $099e2
          39395 => x"7f", -- $099e3
          39396 => x"7f", -- $099e4
          39397 => x"7f", -- $099e5
          39398 => x"7f", -- $099e6
          39399 => x"7f", -- $099e7
          39400 => x"80", -- $099e8
          39401 => x"80", -- $099e9
          39402 => x"80", -- $099ea
          39403 => x"80", -- $099eb
          39404 => x"80", -- $099ec
          39405 => x"80", -- $099ed
          39406 => x"80", -- $099ee
          39407 => x"80", -- $099ef
          39408 => x"80", -- $099f0
          39409 => x"80", -- $099f1
          39410 => x"80", -- $099f2
          39411 => x"80", -- $099f3
          39412 => x"80", -- $099f4
          39413 => x"80", -- $099f5
          39414 => x"80", -- $099f6
          39415 => x"80", -- $099f7
          39416 => x"80", -- $099f8
          39417 => x"7f", -- $099f9
          39418 => x"7f", -- $099fa
          39419 => x"7f", -- $099fb
          39420 => x"7f", -- $099fc
          39421 => x"7f", -- $099fd
          39422 => x"7f", -- $099fe
          39423 => x"7f", -- $099ff
          39424 => x"7f", -- $09a00
          39425 => x"7f", -- $09a01
          39426 => x"7f", -- $09a02
          39427 => x"7f", -- $09a03
          39428 => x"7f", -- $09a04
          39429 => x"7f", -- $09a05
          39430 => x"7f", -- $09a06
          39431 => x"80", -- $09a07
          39432 => x"80", -- $09a08
          39433 => x"80", -- $09a09
          39434 => x"80", -- $09a0a
          39435 => x"80", -- $09a0b
          39436 => x"80", -- $09a0c
          39437 => x"80", -- $09a0d
          39438 => x"80", -- $09a0e
          39439 => x"80", -- $09a0f
          39440 => x"80", -- $09a10
          39441 => x"80", -- $09a11
          39442 => x"80", -- $09a12
          39443 => x"80", -- $09a13
          39444 => x"80", -- $09a14
          39445 => x"80", -- $09a15
          39446 => x"80", -- $09a16
          39447 => x"80", -- $09a17
          39448 => x"80", -- $09a18
          39449 => x"80", -- $09a19
          39450 => x"80", -- $09a1a
          39451 => x"80", -- $09a1b
          39452 => x"80", -- $09a1c
          39453 => x"80", -- $09a1d
          39454 => x"80", -- $09a1e
          39455 => x"80", -- $09a1f
          39456 => x"80", -- $09a20
          39457 => x"80", -- $09a21
          39458 => x"80", -- $09a22
          39459 => x"80", -- $09a23
          39460 => x"80", -- $09a24
          39461 => x"80", -- $09a25
          39462 => x"80", -- $09a26
          39463 => x"80", -- $09a27
          39464 => x"80", -- $09a28
          39465 => x"80", -- $09a29
          39466 => x"80", -- $09a2a
          39467 => x"80", -- $09a2b
          39468 => x"80", -- $09a2c
          39469 => x"80", -- $09a2d
          39470 => x"80", -- $09a2e
          39471 => x"80", -- $09a2f
          39472 => x"80", -- $09a30
          39473 => x"80", -- $09a31
          39474 => x"80", -- $09a32
          39475 => x"80", -- $09a33
          39476 => x"80", -- $09a34
          39477 => x"80", -- $09a35
          39478 => x"80", -- $09a36
          39479 => x"80", -- $09a37
          39480 => x"80", -- $09a38
          39481 => x"80", -- $09a39
          39482 => x"80", -- $09a3a
          39483 => x"80", -- $09a3b
          39484 => x"80", -- $09a3c
          39485 => x"80", -- $09a3d
          39486 => x"80", -- $09a3e
          39487 => x"80", -- $09a3f
          39488 => x"80", -- $09a40
          39489 => x"80", -- $09a41
          39490 => x"80", -- $09a42
          39491 => x"80", -- $09a43
          39492 => x"80", -- $09a44
          39493 => x"80", -- $09a45
          39494 => x"80", -- $09a46
          39495 => x"80", -- $09a47
          39496 => x"80", -- $09a48
          39497 => x"80", -- $09a49
          39498 => x"80", -- $09a4a
          39499 => x"80", -- $09a4b
          39500 => x"80", -- $09a4c
          39501 => x"80", -- $09a4d
          39502 => x"80", -- $09a4e
          39503 => x"80", -- $09a4f
          39504 => x"80", -- $09a50
          39505 => x"80", -- $09a51
          39506 => x"80", -- $09a52
          39507 => x"80", -- $09a53
          39508 => x"80", -- $09a54
          39509 => x"80", -- $09a55
          39510 => x"80", -- $09a56
          39511 => x"80", -- $09a57
          39512 => x"80", -- $09a58
          39513 => x"80", -- $09a59
          39514 => x"80", -- $09a5a
          39515 => x"80", -- $09a5b
          39516 => x"80", -- $09a5c
          39517 => x"80", -- $09a5d
          39518 => x"80", -- $09a5e
          39519 => x"80", -- $09a5f
          39520 => x"80", -- $09a60
          39521 => x"80", -- $09a61
          39522 => x"80", -- $09a62
          39523 => x"80", -- $09a63
          39524 => x"80", -- $09a64
          39525 => x"80", -- $09a65
          39526 => x"80", -- $09a66
          39527 => x"80", -- $09a67
          39528 => x"80", -- $09a68
          39529 => x"80", -- $09a69
          39530 => x"80", -- $09a6a
          39531 => x"80", -- $09a6b
          39532 => x"80", -- $09a6c
          39533 => x"80", -- $09a6d
          39534 => x"80", -- $09a6e
          39535 => x"80", -- $09a6f
          39536 => x"80", -- $09a70
          39537 => x"80", -- $09a71
          39538 => x"80", -- $09a72
          39539 => x"80", -- $09a73
          39540 => x"80", -- $09a74
          39541 => x"80", -- $09a75
          39542 => x"80", -- $09a76
          39543 => x"80", -- $09a77
          39544 => x"80", -- $09a78
          39545 => x"80", -- $09a79
          39546 => x"80", -- $09a7a
          39547 => x"80", -- $09a7b
          39548 => x"80", -- $09a7c
          39549 => x"80", -- $09a7d
          39550 => x"80", -- $09a7e
          39551 => x"80", -- $09a7f
          39552 => x"80", -- $09a80
          39553 => x"80", -- $09a81
          39554 => x"80", -- $09a82
          39555 => x"80", -- $09a83
          39556 => x"80", -- $09a84
          39557 => x"80", -- $09a85
          39558 => x"80", -- $09a86
          39559 => x"80", -- $09a87
          39560 => x"80", -- $09a88
          39561 => x"80", -- $09a89
          39562 => x"80", -- $09a8a
          39563 => x"80", -- $09a8b
          39564 => x"80", -- $09a8c
          39565 => x"80", -- $09a8d
          39566 => x"80", -- $09a8e
          39567 => x"80", -- $09a8f
          39568 => x"80", -- $09a90
          39569 => x"80", -- $09a91
          39570 => x"80", -- $09a92
          39571 => x"80", -- $09a93
          39572 => x"80", -- $09a94
          39573 => x"80", -- $09a95
          39574 => x"80", -- $09a96
          39575 => x"80", -- $09a97
          39576 => x"80", -- $09a98
          39577 => x"80", -- $09a99
          39578 => x"80", -- $09a9a
          39579 => x"80", -- $09a9b
          39580 => x"80", -- $09a9c
          39581 => x"80", -- $09a9d
          39582 => x"80", -- $09a9e
          39583 => x"80", -- $09a9f
          39584 => x"80", -- $09aa0
          39585 => x"80", -- $09aa1
          39586 => x"80", -- $09aa2
          39587 => x"80", -- $09aa3
          39588 => x"80", -- $09aa4
          39589 => x"80", -- $09aa5
          39590 => x"80", -- $09aa6
          39591 => x"80", -- $09aa7
          39592 => x"80", -- $09aa8
          39593 => x"80", -- $09aa9
          39594 => x"80", -- $09aaa
          39595 => x"80", -- $09aab
          39596 => x"80", -- $09aac
          39597 => x"80", -- $09aad
          39598 => x"80", -- $09aae
          39599 => x"80", -- $09aaf
          39600 => x"80", -- $09ab0
          39601 => x"80", -- $09ab1
          39602 => x"80", -- $09ab2
          39603 => x"80", -- $09ab3
          39604 => x"80", -- $09ab4
          39605 => x"80", -- $09ab5
          39606 => x"80", -- $09ab6
          39607 => x"80", -- $09ab7
          39608 => x"80", -- $09ab8
          39609 => x"80", -- $09ab9
          39610 => x"80", -- $09aba
          39611 => x"80", -- $09abb
          39612 => x"80", -- $09abc
          39613 => x"80", -- $09abd
          39614 => x"80", -- $09abe
          39615 => x"80", -- $09abf
          39616 => x"80", -- $09ac0
          39617 => x"80", -- $09ac1
          39618 => x"80", -- $09ac2
          39619 => x"80", -- $09ac3
          39620 => x"80", -- $09ac4
          39621 => x"80", -- $09ac5
          39622 => x"80", -- $09ac6
          39623 => x"80", -- $09ac7
          39624 => x"80", -- $09ac8
          39625 => x"80", -- $09ac9
          39626 => x"80", -- $09aca
          39627 => x"80", -- $09acb
          39628 => x"80", -- $09acc
          39629 => x"80", -- $09acd
          39630 => x"80", -- $09ace
          39631 => x"80", -- $09acf
          39632 => x"80", -- $09ad0
          39633 => x"80", -- $09ad1
          39634 => x"80", -- $09ad2
          39635 => x"80", -- $09ad3
          39636 => x"80", -- $09ad4
          39637 => x"80", -- $09ad5
          39638 => x"80", -- $09ad6
          39639 => x"80", -- $09ad7
          39640 => x"80", -- $09ad8
          39641 => x"80", -- $09ad9
          39642 => x"80", -- $09ada
          39643 => x"80", -- $09adb
          39644 => x"80", -- $09adc
          39645 => x"80", -- $09add
          39646 => x"80", -- $09ade
          39647 => x"80", -- $09adf
          39648 => x"80", -- $09ae0
          39649 => x"80", -- $09ae1
          39650 => x"80", -- $09ae2
          39651 => x"80", -- $09ae3
          39652 => x"80", -- $09ae4
          39653 => x"80", -- $09ae5
          39654 => x"80", -- $09ae6
          39655 => x"80", -- $09ae7
          39656 => x"81", -- $09ae8
          39657 => x"81", -- $09ae9
          39658 => x"81", -- $09aea
          39659 => x"81", -- $09aeb
          39660 => x"81", -- $09aec
          39661 => x"81", -- $09aed
          39662 => x"81", -- $09aee
          39663 => x"81", -- $09aef
          39664 => x"81", -- $09af0
          39665 => x"81", -- $09af1
          39666 => x"81", -- $09af2
          39667 => x"81", -- $09af3
          39668 => x"81", -- $09af4
          39669 => x"81", -- $09af5
          39670 => x"81", -- $09af6
          39671 => x"81", -- $09af7
          39672 => x"81", -- $09af8
          39673 => x"81", -- $09af9
          39674 => x"81", -- $09afa
          39675 => x"81", -- $09afb
          39676 => x"80", -- $09afc
          39677 => x"80", -- $09afd
          39678 => x"80", -- $09afe
          39679 => x"80", -- $09aff
          39680 => x"81", -- $09b00
          39681 => x"81", -- $09b01
          39682 => x"81", -- $09b02
          39683 => x"81", -- $09b03
          39684 => x"81", -- $09b04
          39685 => x"81", -- $09b05
          39686 => x"81", -- $09b06
          39687 => x"81", -- $09b07
          39688 => x"81", -- $09b08
          39689 => x"81", -- $09b09
          39690 => x"81", -- $09b0a
          39691 => x"81", -- $09b0b
          39692 => x"81", -- $09b0c
          39693 => x"81", -- $09b0d
          39694 => x"81", -- $09b0e
          39695 => x"81", -- $09b0f
          39696 => x"81", -- $09b10
          39697 => x"81", -- $09b11
          39698 => x"81", -- $09b12
          39699 => x"81", -- $09b13
          39700 => x"81", -- $09b14
          39701 => x"81", -- $09b15
          39702 => x"81", -- $09b16
          39703 => x"81", -- $09b17
          39704 => x"81", -- $09b18
          39705 => x"81", -- $09b19
          39706 => x"81", -- $09b1a
          39707 => x"81", -- $09b1b
          39708 => x"81", -- $09b1c
          39709 => x"81", -- $09b1d
          39710 => x"81", -- $09b1e
          39711 => x"81", -- $09b1f
          39712 => x"81", -- $09b20
          39713 => x"81", -- $09b21
          39714 => x"80", -- $09b22
          39715 => x"81", -- $09b23
          39716 => x"81", -- $09b24
          39717 => x"81", -- $09b25
          39718 => x"81", -- $09b26
          39719 => x"81", -- $09b27
          39720 => x"81", -- $09b28
          39721 => x"81", -- $09b29
          39722 => x"81", -- $09b2a
          39723 => x"81", -- $09b2b
          39724 => x"81", -- $09b2c
          39725 => x"81", -- $09b2d
          39726 => x"81", -- $09b2e
          39727 => x"81", -- $09b2f
          39728 => x"81", -- $09b30
          39729 => x"81", -- $09b31
          39730 => x"81", -- $09b32
          39731 => x"81", -- $09b33
          39732 => x"81", -- $09b34
          39733 => x"81", -- $09b35
          39734 => x"81", -- $09b36
          39735 => x"81", -- $09b37
          39736 => x"81", -- $09b38
          39737 => x"81", -- $09b39
          39738 => x"81", -- $09b3a
          39739 => x"81", -- $09b3b
          39740 => x"81", -- $09b3c
          39741 => x"81", -- $09b3d
          39742 => x"81", -- $09b3e
          39743 => x"81", -- $09b3f
          39744 => x"81", -- $09b40
          39745 => x"81", -- $09b41
          39746 => x"81", -- $09b42
          39747 => x"81", -- $09b43
          39748 => x"81", -- $09b44
          39749 => x"81", -- $09b45
          39750 => x"81", -- $09b46
          39751 => x"81", -- $09b47
          39752 => x"81", -- $09b48
          39753 => x"81", -- $09b49
          39754 => x"81", -- $09b4a
          39755 => x"81", -- $09b4b
          39756 => x"80", -- $09b4c
          39757 => x"80", -- $09b4d
          39758 => x"80", -- $09b4e
          39759 => x"81", -- $09b4f
          39760 => x"80", -- $09b50
          39761 => x"81", -- $09b51
          39762 => x"81", -- $09b52
          39763 => x"81", -- $09b53
          39764 => x"80", -- $09b54
          39765 => x"81", -- $09b55
          39766 => x"80", -- $09b56
          39767 => x"81", -- $09b57
          39768 => x"81", -- $09b58
          39769 => x"80", -- $09b59
          39770 => x"81", -- $09b5a
          39771 => x"81", -- $09b5b
          39772 => x"80", -- $09b5c
          39773 => x"81", -- $09b5d
          39774 => x"81", -- $09b5e
          39775 => x"81", -- $09b5f
          39776 => x"81", -- $09b60
          39777 => x"81", -- $09b61
          39778 => x"81", -- $09b62
          39779 => x"81", -- $09b63
          39780 => x"80", -- $09b64
          39781 => x"80", -- $09b65
          39782 => x"80", -- $09b66
          39783 => x"80", -- $09b67
          39784 => x"80", -- $09b68
          39785 => x"80", -- $09b69
          39786 => x"80", -- $09b6a
          39787 => x"80", -- $09b6b
          39788 => x"80", -- $09b6c
          39789 => x"80", -- $09b6d
          39790 => x"80", -- $09b6e
          39791 => x"80", -- $09b6f
          39792 => x"80", -- $09b70
          39793 => x"80", -- $09b71
          39794 => x"80", -- $09b72
          39795 => x"80", -- $09b73
          39796 => x"80", -- $09b74
          39797 => x"81", -- $09b75
          39798 => x"81", -- $09b76
          39799 => x"81", -- $09b77
          39800 => x"81", -- $09b78
          39801 => x"81", -- $09b79
          39802 => x"81", -- $09b7a
          39803 => x"81", -- $09b7b
          39804 => x"81", -- $09b7c
          39805 => x"81", -- $09b7d
          39806 => x"81", -- $09b7e
          39807 => x"80", -- $09b7f
          39808 => x"80", -- $09b80
          39809 => x"80", -- $09b81
          39810 => x"80", -- $09b82
          39811 => x"80", -- $09b83
          39812 => x"80", -- $09b84
          39813 => x"80", -- $09b85
          39814 => x"80", -- $09b86
          39815 => x"80", -- $09b87
          39816 => x"80", -- $09b88
          39817 => x"80", -- $09b89
          39818 => x"80", -- $09b8a
          39819 => x"80", -- $09b8b
          39820 => x"80", -- $09b8c
          39821 => x"80", -- $09b8d
          39822 => x"80", -- $09b8e
          39823 => x"80", -- $09b8f
          39824 => x"80", -- $09b90
          39825 => x"80", -- $09b91
          39826 => x"80", -- $09b92
          39827 => x"80", -- $09b93
          39828 => x"80", -- $09b94
          39829 => x"80", -- $09b95
          39830 => x"80", -- $09b96
          39831 => x"80", -- $09b97
          39832 => x"80", -- $09b98
          39833 => x"80", -- $09b99
          39834 => x"80", -- $09b9a
          39835 => x"80", -- $09b9b
          39836 => x"80", -- $09b9c
          39837 => x"80", -- $09b9d
          39838 => x"80", -- $09b9e
          39839 => x"80", -- $09b9f
          39840 => x"80", -- $09ba0
          39841 => x"80", -- $09ba1
          39842 => x"80", -- $09ba2
          39843 => x"80", -- $09ba3
          39844 => x"80", -- $09ba4
          39845 => x"80", -- $09ba5
          39846 => x"80", -- $09ba6
          39847 => x"80", -- $09ba7
          39848 => x"80", -- $09ba8
          39849 => x"80", -- $09ba9
          39850 => x"80", -- $09baa
          39851 => x"80", -- $09bab
          39852 => x"80", -- $09bac
          39853 => x"80", -- $09bad
          39854 => x"80", -- $09bae
          39855 => x"80", -- $09baf
          39856 => x"80", -- $09bb0
          39857 => x"80", -- $09bb1
          39858 => x"80", -- $09bb2
          39859 => x"80", -- $09bb3
          39860 => x"80", -- $09bb4
          39861 => x"80", -- $09bb5
          39862 => x"80", -- $09bb6
          39863 => x"80", -- $09bb7
          39864 => x"80", -- $09bb8
          39865 => x"80", -- $09bb9
          39866 => x"80", -- $09bba
          39867 => x"80", -- $09bbb
          39868 => x"80", -- $09bbc
          39869 => x"80", -- $09bbd
          39870 => x"80", -- $09bbe
          39871 => x"80", -- $09bbf
          39872 => x"80", -- $09bc0
          39873 => x"80", -- $09bc1
          39874 => x"80", -- $09bc2
          39875 => x"80", -- $09bc3
          39876 => x"80", -- $09bc4
          39877 => x"80", -- $09bc5
          39878 => x"80", -- $09bc6
          39879 => x"80", -- $09bc7
          39880 => x"80", -- $09bc8
          39881 => x"80", -- $09bc9
          39882 => x"80", -- $09bca
          39883 => x"80", -- $09bcb
          39884 => x"80", -- $09bcc
          39885 => x"80", -- $09bcd
          39886 => x"80", -- $09bce
          39887 => x"80", -- $09bcf
          39888 => x"80", -- $09bd0
          39889 => x"80", -- $09bd1
          39890 => x"80", -- $09bd2
          39891 => x"80", -- $09bd3
          39892 => x"80", -- $09bd4
          39893 => x"80", -- $09bd5
          39894 => x"80", -- $09bd6
          39895 => x"80", -- $09bd7
          39896 => x"80", -- $09bd8
          39897 => x"80", -- $09bd9
          39898 => x"80", -- $09bda
          39899 => x"80", -- $09bdb
          39900 => x"80", -- $09bdc
          39901 => x"80", -- $09bdd
          39902 => x"80", -- $09bde
          39903 => x"80", -- $09bdf
          39904 => x"80", -- $09be0
          39905 => x"80", -- $09be1
          39906 => x"80", -- $09be2
          39907 => x"80", -- $09be3
          39908 => x"80", -- $09be4
          39909 => x"80", -- $09be5
          39910 => x"80", -- $09be6
          39911 => x"80", -- $09be7
          39912 => x"80", -- $09be8
          39913 => x"80", -- $09be9
          39914 => x"80", -- $09bea
          39915 => x"80", -- $09beb
          39916 => x"80", -- $09bec
          39917 => x"80", -- $09bed
          39918 => x"80", -- $09bee
          39919 => x"80", -- $09bef
          39920 => x"7f", -- $09bf0
          39921 => x"80", -- $09bf1
          39922 => x"80", -- $09bf2
          39923 => x"80", -- $09bf3
          39924 => x"80", -- $09bf4
          39925 => x"80", -- $09bf5
          39926 => x"80", -- $09bf6
          39927 => x"80", -- $09bf7
          39928 => x"80", -- $09bf8
          39929 => x"80", -- $09bf9
          39930 => x"80", -- $09bfa
          39931 => x"80", -- $09bfb
          39932 => x"80", -- $09bfc
          39933 => x"80", -- $09bfd
          39934 => x"80", -- $09bfe
          39935 => x"80", -- $09bff
          39936 => x"80", -- $09c00
          39937 => x"80", -- $09c01
          39938 => x"80", -- $09c02
          39939 => x"80", -- $09c03
          39940 => x"80", -- $09c04
          39941 => x"80", -- $09c05
          39942 => x"80", -- $09c06
          39943 => x"80", -- $09c07
          39944 => x"80", -- $09c08
          39945 => x"80", -- $09c09
          39946 => x"80", -- $09c0a
          39947 => x"7f", -- $09c0b
          39948 => x"7f", -- $09c0c
          39949 => x"80", -- $09c0d
          39950 => x"80", -- $09c0e
          39951 => x"80", -- $09c0f
          39952 => x"80", -- $09c10
          39953 => x"80", -- $09c11
          39954 => x"80", -- $09c12
          39955 => x"80", -- $09c13
          39956 => x"80", -- $09c14
          39957 => x"80", -- $09c15
          39958 => x"80", -- $09c16
          39959 => x"80", -- $09c17
          39960 => x"80", -- $09c18
          39961 => x"80", -- $09c19
          39962 => x"80", -- $09c1a
          39963 => x"80", -- $09c1b
          39964 => x"80", -- $09c1c
          39965 => x"80", -- $09c1d
          39966 => x"80", -- $09c1e
          39967 => x"80", -- $09c1f
          39968 => x"80", -- $09c20
          39969 => x"80", -- $09c21
          39970 => x"80", -- $09c22
          39971 => x"80", -- $09c23
          39972 => x"80", -- $09c24
          39973 => x"7f", -- $09c25
          39974 => x"7f", -- $09c26
          39975 => x"7f", -- $09c27
          39976 => x"7f", -- $09c28
          39977 => x"7f", -- $09c29
          39978 => x"7f", -- $09c2a
          39979 => x"7f", -- $09c2b
          39980 => x"7f", -- $09c2c
          39981 => x"80", -- $09c2d
          39982 => x"80", -- $09c2e
          39983 => x"80", -- $09c2f
          39984 => x"80", -- $09c30
          39985 => x"80", -- $09c31
          39986 => x"80", -- $09c32
          39987 => x"80", -- $09c33
          39988 => x"80", -- $09c34
          39989 => x"80", -- $09c35
          39990 => x"80", -- $09c36
          39991 => x"80", -- $09c37
          39992 => x"80", -- $09c38
          39993 => x"80", -- $09c39
          39994 => x"80", -- $09c3a
          39995 => x"80", -- $09c3b
          39996 => x"80", -- $09c3c
          39997 => x"80", -- $09c3d
          39998 => x"7f", -- $09c3e
          39999 => x"7f", -- $09c3f
          40000 => x"7f", -- $09c40
          40001 => x"7f", -- $09c41
          40002 => x"7f", -- $09c42
          40003 => x"7f", -- $09c43
          40004 => x"7f", -- $09c44
          40005 => x"7f", -- $09c45
          40006 => x"7f", -- $09c46
          40007 => x"7f", -- $09c47
          40008 => x"7f", -- $09c48
          40009 => x"7f", -- $09c49
          40010 => x"7f", -- $09c4a
          40011 => x"7f", -- $09c4b
          40012 => x"7f", -- $09c4c
          40013 => x"7f", -- $09c4d
          40014 => x"7f", -- $09c4e
          40015 => x"7f", -- $09c4f
          40016 => x"7f", -- $09c50
          40017 => x"7f", -- $09c51
          40018 => x"7f", -- $09c52
          40019 => x"7f", -- $09c53
          40020 => x"7f", -- $09c54
          40021 => x"7f", -- $09c55
          40022 => x"7f", -- $09c56
          40023 => x"7f", -- $09c57
          40024 => x"7f", -- $09c58
          40025 => x"7f", -- $09c59
          40026 => x"7f", -- $09c5a
          40027 => x"7e", -- $09c5b
          40028 => x"7e", -- $09c5c
          40029 => x"7e", -- $09c5d
          40030 => x"7e", -- $09c5e
          40031 => x"7e", -- $09c5f
          40032 => x"7f", -- $09c60
          40033 => x"7f", -- $09c61
          40034 => x"7f", -- $09c62
          40035 => x"7f", -- $09c63
          40036 => x"7f", -- $09c64
          40037 => x"7f", -- $09c65
          40038 => x"7f", -- $09c66
          40039 => x"7f", -- $09c67
          40040 => x"7f", -- $09c68
          40041 => x"7f", -- $09c69
          40042 => x"7f", -- $09c6a
          40043 => x"7f", -- $09c6b
          40044 => x"7f", -- $09c6c
          40045 => x"7f", -- $09c6d
          40046 => x"7f", -- $09c6e
          40047 => x"7f", -- $09c6f
          40048 => x"7f", -- $09c70
          40049 => x"7f", -- $09c71
          40050 => x"7f", -- $09c72
          40051 => x"7f", -- $09c73
          40052 => x"7f", -- $09c74
          40053 => x"7f", -- $09c75
          40054 => x"7f", -- $09c76
          40055 => x"7e", -- $09c77
          40056 => x"7e", -- $09c78
          40057 => x"7e", -- $09c79
          40058 => x"7f", -- $09c7a
          40059 => x"7f", -- $09c7b
          40060 => x"7f", -- $09c7c
          40061 => x"7f", -- $09c7d
          40062 => x"7f", -- $09c7e
          40063 => x"7f", -- $09c7f
          40064 => x"7f", -- $09c80
          40065 => x"7f", -- $09c81
          40066 => x"7f", -- $09c82
          40067 => x"7f", -- $09c83
          40068 => x"7f", -- $09c84
          40069 => x"7f", -- $09c85
          40070 => x"7f", -- $09c86
          40071 => x"7f", -- $09c87
          40072 => x"7f", -- $09c88
          40073 => x"7f", -- $09c89
          40074 => x"7f", -- $09c8a
          40075 => x"7f", -- $09c8b
          40076 => x"7f", -- $09c8c
          40077 => x"7f", -- $09c8d
          40078 => x"7f", -- $09c8e
          40079 => x"7f", -- $09c8f
          40080 => x"7f", -- $09c90
          40081 => x"7f", -- $09c91
          40082 => x"7f", -- $09c92
          40083 => x"7e", -- $09c93
          40084 => x"7f", -- $09c94
          40085 => x"7f", -- $09c95
          40086 => x"7f", -- $09c96
          40087 => x"7f", -- $09c97
          40088 => x"7f", -- $09c98
          40089 => x"7f", -- $09c99
          40090 => x"7f", -- $09c9a
          40091 => x"7f", -- $09c9b
          40092 => x"7f", -- $09c9c
          40093 => x"7f", -- $09c9d
          40094 => x"7f", -- $09c9e
          40095 => x"7f", -- $09c9f
          40096 => x"80", -- $09ca0
          40097 => x"80", -- $09ca1
          40098 => x"80", -- $09ca2
          40099 => x"80", -- $09ca3
          40100 => x"80", -- $09ca4
          40101 => x"80", -- $09ca5
          40102 => x"80", -- $09ca6
          40103 => x"80", -- $09ca7
          40104 => x"80", -- $09ca8
          40105 => x"80", -- $09ca9
          40106 => x"80", -- $09caa
          40107 => x"7f", -- $09cab
          40108 => x"7f", -- $09cac
          40109 => x"7f", -- $09cad
          40110 => x"7f", -- $09cae
          40111 => x"7f", -- $09caf
          40112 => x"7f", -- $09cb0
          40113 => x"7f", -- $09cb1
          40114 => x"7f", -- $09cb2
          40115 => x"7f", -- $09cb3
          40116 => x"7f", -- $09cb4
          40117 => x"80", -- $09cb5
          40118 => x"80", -- $09cb6
          40119 => x"80", -- $09cb7
          40120 => x"80", -- $09cb8
          40121 => x"80", -- $09cb9
          40122 => x"80", -- $09cba
          40123 => x"80", -- $09cbb
          40124 => x"80", -- $09cbc
          40125 => x"80", -- $09cbd
          40126 => x"80", -- $09cbe
          40127 => x"80", -- $09cbf
          40128 => x"80", -- $09cc0
          40129 => x"80", -- $09cc1
          40130 => x"80", -- $09cc2
          40131 => x"80", -- $09cc3
          40132 => x"80", -- $09cc4
          40133 => x"80", -- $09cc5
          40134 => x"80", -- $09cc6
          40135 => x"7f", -- $09cc7
          40136 => x"80", -- $09cc8
          40137 => x"80", -- $09cc9
          40138 => x"80", -- $09cca
          40139 => x"80", -- $09ccb
          40140 => x"80", -- $09ccc
          40141 => x"80", -- $09ccd
          40142 => x"80", -- $09cce
          40143 => x"80", -- $09ccf
          40144 => x"80", -- $09cd0
          40145 => x"80", -- $09cd1
          40146 => x"80", -- $09cd2
          40147 => x"80", -- $09cd3
          40148 => x"80", -- $09cd4
          40149 => x"80", -- $09cd5
          40150 => x"80", -- $09cd6
          40151 => x"80", -- $09cd7
          40152 => x"80", -- $09cd8
          40153 => x"80", -- $09cd9
          40154 => x"80", -- $09cda
          40155 => x"80", -- $09cdb
          40156 => x"80", -- $09cdc
          40157 => x"80", -- $09cdd
          40158 => x"80", -- $09cde
          40159 => x"80", -- $09cdf
          40160 => x"80", -- $09ce0
          40161 => x"80", -- $09ce1
          40162 => x"80", -- $09ce2
          40163 => x"80", -- $09ce3
          40164 => x"80", -- $09ce4
          40165 => x"80", -- $09ce5
          40166 => x"80", -- $09ce6
          40167 => x"80", -- $09ce7
          40168 => x"80", -- $09ce8
          40169 => x"80", -- $09ce9
          40170 => x"80", -- $09cea
          40171 => x"80", -- $09ceb
          40172 => x"80", -- $09cec
          40173 => x"80", -- $09ced
          40174 => x"80", -- $09cee
          40175 => x"80", -- $09cef
          40176 => x"80", -- $09cf0
          40177 => x"80", -- $09cf1
          40178 => x"80", -- $09cf2
          40179 => x"80", -- $09cf3
          40180 => x"80", -- $09cf4
          40181 => x"80", -- $09cf5
          40182 => x"80", -- $09cf6
          40183 => x"80", -- $09cf7
          40184 => x"80", -- $09cf8
          40185 => x"80", -- $09cf9
          40186 => x"80", -- $09cfa
          40187 => x"80", -- $09cfb
          40188 => x"80", -- $09cfc
          40189 => x"80", -- $09cfd
          40190 => x"80", -- $09cfe
          40191 => x"80", -- $09cff
          40192 => x"80", -- $09d00
          40193 => x"80", -- $09d01
          40194 => x"80", -- $09d02
          40195 => x"80", -- $09d03
          40196 => x"7f", -- $09d04
          40197 => x"7f", -- $09d05
          40198 => x"7f", -- $09d06
          40199 => x"7f", -- $09d07
          40200 => x"7f", -- $09d08
          40201 => x"7f", -- $09d09
          40202 => x"80", -- $09d0a
          40203 => x"80", -- $09d0b
          40204 => x"80", -- $09d0c
          40205 => x"80", -- $09d0d
          40206 => x"80", -- $09d0e
          40207 => x"80", -- $09d0f
          40208 => x"80", -- $09d10
          40209 => x"80", -- $09d11
          40210 => x"80", -- $09d12
          40211 => x"80", -- $09d13
          40212 => x"80", -- $09d14
          40213 => x"80", -- $09d15
          40214 => x"80", -- $09d16
          40215 => x"7f", -- $09d17
          40216 => x"80", -- $09d18
          40217 => x"80", -- $09d19
          40218 => x"80", -- $09d1a
          40219 => x"80", -- $09d1b
          40220 => x"80", -- $09d1c
          40221 => x"80", -- $09d1d
          40222 => x"7f", -- $09d1e
          40223 => x"80", -- $09d1f
          40224 => x"80", -- $09d20
          40225 => x"7f", -- $09d21
          40226 => x"80", -- $09d22
          40227 => x"80", -- $09d23
          40228 => x"7f", -- $09d24
          40229 => x"80", -- $09d25
          40230 => x"80", -- $09d26
          40231 => x"80", -- $09d27
          40232 => x"80", -- $09d28
          40233 => x"80", -- $09d29
          40234 => x"80", -- $09d2a
          40235 => x"80", -- $09d2b
          40236 => x"80", -- $09d2c
          40237 => x"80", -- $09d2d
          40238 => x"80", -- $09d2e
          40239 => x"80", -- $09d2f
          40240 => x"80", -- $09d30
          40241 => x"80", -- $09d31
          40242 => x"80", -- $09d32
          40243 => x"80", -- $09d33
          40244 => x"80", -- $09d34
          40245 => x"80", -- $09d35
          40246 => x"80", -- $09d36
          40247 => x"80", -- $09d37
          40248 => x"80", -- $09d38
          40249 => x"80", -- $09d39
          40250 => x"80", -- $09d3a
          40251 => x"80", -- $09d3b
          40252 => x"80", -- $09d3c
          40253 => x"80", -- $09d3d
          40254 => x"80", -- $09d3e
          40255 => x"80", -- $09d3f
          40256 => x"80", -- $09d40
          40257 => x"80", -- $09d41
          40258 => x"80", -- $09d42
          40259 => x"80", -- $09d43
          40260 => x"80", -- $09d44
          40261 => x"80", -- $09d45
          40262 => x"80", -- $09d46
          40263 => x"80", -- $09d47
          40264 => x"80", -- $09d48
          40265 => x"80", -- $09d49
          40266 => x"80", -- $09d4a
          40267 => x"80", -- $09d4b
          40268 => x"80", -- $09d4c
          40269 => x"80", -- $09d4d
          40270 => x"80", -- $09d4e
          40271 => x"80", -- $09d4f
          40272 => x"80", -- $09d50
          40273 => x"80", -- $09d51
          40274 => x"80", -- $09d52
          40275 => x"80", -- $09d53
          40276 => x"80", -- $09d54
          40277 => x"80", -- $09d55
          40278 => x"80", -- $09d56
          40279 => x"80", -- $09d57
          40280 => x"80", -- $09d58
          40281 => x"80", -- $09d59
          40282 => x"80", -- $09d5a
          40283 => x"80", -- $09d5b
          40284 => x"80", -- $09d5c
          40285 => x"80", -- $09d5d
          40286 => x"80", -- $09d5e
          40287 => x"80", -- $09d5f
          40288 => x"80", -- $09d60
          40289 => x"80", -- $09d61
          40290 => x"80", -- $09d62
          40291 => x"80", -- $09d63
          40292 => x"80", -- $09d64
          40293 => x"80", -- $09d65
          40294 => x"80", -- $09d66
          40295 => x"80", -- $09d67
          40296 => x"80", -- $09d68
          40297 => x"80", -- $09d69
          40298 => x"80", -- $09d6a
          40299 => x"80", -- $09d6b
          40300 => x"80", -- $09d6c
          40301 => x"80", -- $09d6d
          40302 => x"80", -- $09d6e
          40303 => x"81", -- $09d6f
          40304 => x"81", -- $09d70
          40305 => x"81", -- $09d71
          40306 => x"81", -- $09d72
          40307 => x"80", -- $09d73
          40308 => x"81", -- $09d74
          40309 => x"81", -- $09d75
          40310 => x"80", -- $09d76
          40311 => x"81", -- $09d77
          40312 => x"81", -- $09d78
          40313 => x"81", -- $09d79
          40314 => x"81", -- $09d7a
          40315 => x"81", -- $09d7b
          40316 => x"80", -- $09d7c
          40317 => x"81", -- $09d7d
          40318 => x"81", -- $09d7e
          40319 => x"81", -- $09d7f
          40320 => x"81", -- $09d80
          40321 => x"81", -- $09d81
          40322 => x"81", -- $09d82
          40323 => x"81", -- $09d83
          40324 => x"81", -- $09d84
          40325 => x"81", -- $09d85
          40326 => x"81", -- $09d86
          40327 => x"81", -- $09d87
          40328 => x"81", -- $09d88
          40329 => x"81", -- $09d89
          40330 => x"81", -- $09d8a
          40331 => x"81", -- $09d8b
          40332 => x"81", -- $09d8c
          40333 => x"81", -- $09d8d
          40334 => x"81", -- $09d8e
          40335 => x"81", -- $09d8f
          40336 => x"81", -- $09d90
          40337 => x"81", -- $09d91
          40338 => x"81", -- $09d92
          40339 => x"81", -- $09d93
          40340 => x"81", -- $09d94
          40341 => x"81", -- $09d95
          40342 => x"81", -- $09d96
          40343 => x"81", -- $09d97
          40344 => x"81", -- $09d98
          40345 => x"81", -- $09d99
          40346 => x"81", -- $09d9a
          40347 => x"81", -- $09d9b
          40348 => x"81", -- $09d9c
          40349 => x"81", -- $09d9d
          40350 => x"81", -- $09d9e
          40351 => x"81", -- $09d9f
          40352 => x"81", -- $09da0
          40353 => x"81", -- $09da1
          40354 => x"81", -- $09da2
          40355 => x"81", -- $09da3
          40356 => x"81", -- $09da4
          40357 => x"81", -- $09da5
          40358 => x"81", -- $09da6
          40359 => x"81", -- $09da7
          40360 => x"81", -- $09da8
          40361 => x"81", -- $09da9
          40362 => x"81", -- $09daa
          40363 => x"81", -- $09dab
          40364 => x"81", -- $09dac
          40365 => x"81", -- $09dad
          40366 => x"81", -- $09dae
          40367 => x"81", -- $09daf
          40368 => x"80", -- $09db0
          40369 => x"80", -- $09db1
          40370 => x"81", -- $09db2
          40371 => x"80", -- $09db3
          40372 => x"80", -- $09db4
          40373 => x"81", -- $09db5
          40374 => x"81", -- $09db6
          40375 => x"81", -- $09db7
          40376 => x"81", -- $09db8
          40377 => x"81", -- $09db9
          40378 => x"81", -- $09dba
          40379 => x"81", -- $09dbb
          40380 => x"81", -- $09dbc
          40381 => x"81", -- $09dbd
          40382 => x"81", -- $09dbe
          40383 => x"81", -- $09dbf
          40384 => x"81", -- $09dc0
          40385 => x"81", -- $09dc1
          40386 => x"81", -- $09dc2
          40387 => x"81", -- $09dc3
          40388 => x"81", -- $09dc4
          40389 => x"81", -- $09dc5
          40390 => x"81", -- $09dc6
          40391 => x"81", -- $09dc7
          40392 => x"81", -- $09dc8
          40393 => x"81", -- $09dc9
          40394 => x"81", -- $09dca
          40395 => x"81", -- $09dcb
          40396 => x"80", -- $09dcc
          40397 => x"81", -- $09dcd
          40398 => x"80", -- $09dce
          40399 => x"81", -- $09dcf
          40400 => x"81", -- $09dd0
          40401 => x"81", -- $09dd1
          40402 => x"81", -- $09dd2
          40403 => x"81", -- $09dd3
          40404 => x"81", -- $09dd4
          40405 => x"81", -- $09dd5
          40406 => x"81", -- $09dd6
          40407 => x"81", -- $09dd7
          40408 => x"81", -- $09dd8
          40409 => x"81", -- $09dd9
          40410 => x"81", -- $09dda
          40411 => x"81", -- $09ddb
          40412 => x"81", -- $09ddc
          40413 => x"81", -- $09ddd
          40414 => x"81", -- $09dde
          40415 => x"81", -- $09ddf
          40416 => x"81", -- $09de0
          40417 => x"81", -- $09de1
          40418 => x"81", -- $09de2
          40419 => x"81", -- $09de3
          40420 => x"81", -- $09de4
          40421 => x"81", -- $09de5
          40422 => x"81", -- $09de6
          40423 => x"80", -- $09de7
          40424 => x"81", -- $09de8
          40425 => x"80", -- $09de9
          40426 => x"80", -- $09dea
          40427 => x"81", -- $09deb
          40428 => x"81", -- $09dec
          40429 => x"81", -- $09ded
          40430 => x"81", -- $09dee
          40431 => x"81", -- $09def
          40432 => x"81", -- $09df0
          40433 => x"81", -- $09df1
          40434 => x"81", -- $09df2
          40435 => x"81", -- $09df3
          40436 => x"81", -- $09df4
          40437 => x"81", -- $09df5
          40438 => x"81", -- $09df6
          40439 => x"81", -- $09df7
          40440 => x"81", -- $09df8
          40441 => x"81", -- $09df9
          40442 => x"81", -- $09dfa
          40443 => x"81", -- $09dfb
          40444 => x"81", -- $09dfc
          40445 => x"81", -- $09dfd
          40446 => x"81", -- $09dfe
          40447 => x"81", -- $09dff
          40448 => x"81", -- $09e00
          40449 => x"81", -- $09e01
          40450 => x"81", -- $09e02
          40451 => x"81", -- $09e03
          40452 => x"81", -- $09e04
          40453 => x"81", -- $09e05
          40454 => x"81", -- $09e06
          40455 => x"81", -- $09e07
          40456 => x"81", -- $09e08
          40457 => x"81", -- $09e09
          40458 => x"81", -- $09e0a
          40459 => x"80", -- $09e0b
          40460 => x"81", -- $09e0c
          40461 => x"81", -- $09e0d
          40462 => x"81", -- $09e0e
          40463 => x"81", -- $09e0f
          40464 => x"81", -- $09e10
          40465 => x"81", -- $09e11
          40466 => x"81", -- $09e12
          40467 => x"81", -- $09e13
          40468 => x"81", -- $09e14
          40469 => x"81", -- $09e15
          40470 => x"81", -- $09e16
          40471 => x"81", -- $09e17
          40472 => x"81", -- $09e18
          40473 => x"81", -- $09e19
          40474 => x"81", -- $09e1a
          40475 => x"80", -- $09e1b
          40476 => x"80", -- $09e1c
          40477 => x"80", -- $09e1d
          40478 => x"80", -- $09e1e
          40479 => x"80", -- $09e1f
          40480 => x"80", -- $09e20
          40481 => x"80", -- $09e21
          40482 => x"80", -- $09e22
          40483 => x"80", -- $09e23
          40484 => x"80", -- $09e24
          40485 => x"80", -- $09e25
          40486 => x"80", -- $09e26
          40487 => x"80", -- $09e27
          40488 => x"80", -- $09e28
          40489 => x"81", -- $09e29
          40490 => x"81", -- $09e2a
          40491 => x"81", -- $09e2b
          40492 => x"81", -- $09e2c
          40493 => x"81", -- $09e2d
          40494 => x"81", -- $09e2e
          40495 => x"81", -- $09e2f
          40496 => x"81", -- $09e30
          40497 => x"81", -- $09e31
          40498 => x"80", -- $09e32
          40499 => x"81", -- $09e33
          40500 => x"81", -- $09e34
          40501 => x"81", -- $09e35
          40502 => x"81", -- $09e36
          40503 => x"81", -- $09e37
          40504 => x"81", -- $09e38
          40505 => x"81", -- $09e39
          40506 => x"80", -- $09e3a
          40507 => x"80", -- $09e3b
          40508 => x"80", -- $09e3c
          40509 => x"80", -- $09e3d
          40510 => x"80", -- $09e3e
          40511 => x"80", -- $09e3f
          40512 => x"80", -- $09e40
          40513 => x"80", -- $09e41
          40514 => x"81", -- $09e42
          40515 => x"81", -- $09e43
          40516 => x"81", -- $09e44
          40517 => x"81", -- $09e45
          40518 => x"81", -- $09e46
          40519 => x"81", -- $09e47
          40520 => x"81", -- $09e48
          40521 => x"81", -- $09e49
          40522 => x"81", -- $09e4a
          40523 => x"81", -- $09e4b
          40524 => x"81", -- $09e4c
          40525 => x"81", -- $09e4d
          40526 => x"81", -- $09e4e
          40527 => x"81", -- $09e4f
          40528 => x"81", -- $09e50
          40529 => x"81", -- $09e51
          40530 => x"81", -- $09e52
          40531 => x"81", -- $09e53
          40532 => x"81", -- $09e54
          40533 => x"81", -- $09e55
          40534 => x"81", -- $09e56
          40535 => x"81", -- $09e57
          40536 => x"80", -- $09e58
          40537 => x"80", -- $09e59
          40538 => x"80", -- $09e5a
          40539 => x"80", -- $09e5b
          40540 => x"80", -- $09e5c
          40541 => x"80", -- $09e5d
          40542 => x"81", -- $09e5e
          40543 => x"81", -- $09e5f
          40544 => x"81", -- $09e60
          40545 => x"81", -- $09e61
          40546 => x"81", -- $09e62
          40547 => x"81", -- $09e63
          40548 => x"81", -- $09e64
          40549 => x"81", -- $09e65
          40550 => x"81", -- $09e66
          40551 => x"81", -- $09e67
          40552 => x"81", -- $09e68
          40553 => x"81", -- $09e69
          40554 => x"81", -- $09e6a
          40555 => x"81", -- $09e6b
          40556 => x"81", -- $09e6c
          40557 => x"81", -- $09e6d
          40558 => x"81", -- $09e6e
          40559 => x"81", -- $09e6f
          40560 => x"81", -- $09e70
          40561 => x"80", -- $09e71
          40562 => x"80", -- $09e72
          40563 => x"80", -- $09e73
          40564 => x"80", -- $09e74
          40565 => x"80", -- $09e75
          40566 => x"80", -- $09e76
          40567 => x"80", -- $09e77
          40568 => x"80", -- $09e78
          40569 => x"80", -- $09e79
          40570 => x"80", -- $09e7a
          40571 => x"80", -- $09e7b
          40572 => x"81", -- $09e7c
          40573 => x"81", -- $09e7d
          40574 => x"80", -- $09e7e
          40575 => x"81", -- $09e7f
          40576 => x"81", -- $09e80
          40577 => x"80", -- $09e81
          40578 => x"80", -- $09e82
          40579 => x"80", -- $09e83
          40580 => x"80", -- $09e84
          40581 => x"80", -- $09e85
          40582 => x"80", -- $09e86
          40583 => x"80", -- $09e87
          40584 => x"80", -- $09e88
          40585 => x"80", -- $09e89
          40586 => x"80", -- $09e8a
          40587 => x"80", -- $09e8b
          40588 => x"80", -- $09e8c
          40589 => x"80", -- $09e8d
          40590 => x"80", -- $09e8e
          40591 => x"80", -- $09e8f
          40592 => x"80", -- $09e90
          40593 => x"80", -- $09e91
          40594 => x"80", -- $09e92
          40595 => x"80", -- $09e93
          40596 => x"80", -- $09e94
          40597 => x"80", -- $09e95
          40598 => x"80", -- $09e96
          40599 => x"80", -- $09e97
          40600 => x"80", -- $09e98
          40601 => x"80", -- $09e99
          40602 => x"80", -- $09e9a
          40603 => x"80", -- $09e9b
          40604 => x"80", -- $09e9c
          40605 => x"80", -- $09e9d
          40606 => x"80", -- $09e9e
          40607 => x"80", -- $09e9f
          40608 => x"80", -- $09ea0
          40609 => x"80", -- $09ea1
          40610 => x"80", -- $09ea2
          40611 => x"80", -- $09ea3
          40612 => x"80", -- $09ea4
          40613 => x"80", -- $09ea5
          40614 => x"80", -- $09ea6
          40615 => x"80", -- $09ea7
          40616 => x"80", -- $09ea8
          40617 => x"80", -- $09ea9
          40618 => x"80", -- $09eaa
          40619 => x"80", -- $09eab
          40620 => x"80", -- $09eac
          40621 => x"80", -- $09ead
          40622 => x"80", -- $09eae
          40623 => x"80", -- $09eaf
          40624 => x"7f", -- $09eb0
          40625 => x"7f", -- $09eb1
          40626 => x"7f", -- $09eb2
          40627 => x"7f", -- $09eb3
          40628 => x"7f", -- $09eb4
          40629 => x"7f", -- $09eb5
          40630 => x"7f", -- $09eb6
          40631 => x"7f", -- $09eb7
          40632 => x"7f", -- $09eb8
          40633 => x"7f", -- $09eb9
          40634 => x"80", -- $09eba
          40635 => x"80", -- $09ebb
          40636 => x"7f", -- $09ebc
          40637 => x"7f", -- $09ebd
          40638 => x"7f", -- $09ebe
          40639 => x"7f", -- $09ebf
          40640 => x"7f", -- $09ec0
          40641 => x"7f", -- $09ec1
          40642 => x"7f", -- $09ec2
          40643 => x"7f", -- $09ec3
          40644 => x"7f", -- $09ec4
          40645 => x"7f", -- $09ec5
          40646 => x"7f", -- $09ec6
          40647 => x"7f", -- $09ec7
          40648 => x"7f", -- $09ec8
          40649 => x"7f", -- $09ec9
          40650 => x"7f", -- $09eca
          40651 => x"7f", -- $09ecb
          40652 => x"7f", -- $09ecc
          40653 => x"7f", -- $09ecd
          40654 => x"7f", -- $09ece
          40655 => x"7f", -- $09ecf
          40656 => x"7f", -- $09ed0
          40657 => x"7f", -- $09ed1
          40658 => x"7f", -- $09ed2
          40659 => x"7f", -- $09ed3
          40660 => x"7f", -- $09ed4
          40661 => x"7f", -- $09ed5
          40662 => x"7f", -- $09ed6
          40663 => x"7f", -- $09ed7
          40664 => x"7f", -- $09ed8
          40665 => x"7f", -- $09ed9
          40666 => x"7f", -- $09eda
          40667 => x"7f", -- $09edb
          40668 => x"7f", -- $09edc
          40669 => x"7f", -- $09edd
          40670 => x"7f", -- $09ede
          40671 => x"7f", -- $09edf
          40672 => x"7f", -- $09ee0
          40673 => x"7f", -- $09ee1
          40674 => x"7f", -- $09ee2
          40675 => x"7f", -- $09ee3
          40676 => x"7f", -- $09ee4
          40677 => x"7f", -- $09ee5
          40678 => x"7f", -- $09ee6
          40679 => x"7f", -- $09ee7
          40680 => x"7f", -- $09ee8
          40681 => x"7f", -- $09ee9
          40682 => x"7f", -- $09eea
          40683 => x"7f", -- $09eeb
          40684 => x"7f", -- $09eec
          40685 => x"7f", -- $09eed
          40686 => x"7f", -- $09eee
          40687 => x"7f", -- $09eef
          40688 => x"7f", -- $09ef0
          40689 => x"7f", -- $09ef1
          40690 => x"7f", -- $09ef2
          40691 => x"7f", -- $09ef3
          40692 => x"7f", -- $09ef4
          40693 => x"7f", -- $09ef5
          40694 => x"7f", -- $09ef6
          40695 => x"7f", -- $09ef7
          40696 => x"7f", -- $09ef8
          40697 => x"7f", -- $09ef9
          40698 => x"7f", -- $09efa
          40699 => x"7f", -- $09efb
          40700 => x"7f", -- $09efc
          40701 => x"7f", -- $09efd
          40702 => x"7f", -- $09efe
          40703 => x"7f", -- $09eff
          40704 => x"7f", -- $09f00
          40705 => x"7f", -- $09f01
          40706 => x"7f", -- $09f02
          40707 => x"7f", -- $09f03
          40708 => x"7f", -- $09f04
          40709 => x"7f", -- $09f05
          40710 => x"7f", -- $09f06
          40711 => x"7f", -- $09f07
          40712 => x"7f", -- $09f08
          40713 => x"7f", -- $09f09
          40714 => x"7f", -- $09f0a
          40715 => x"7f", -- $09f0b
          40716 => x"7f", -- $09f0c
          40717 => x"7f", -- $09f0d
          40718 => x"7f", -- $09f0e
          40719 => x"7f", -- $09f0f
          40720 => x"7f", -- $09f10
          40721 => x"7f", -- $09f11
          40722 => x"7f", -- $09f12
          40723 => x"7f", -- $09f13
          40724 => x"7f", -- $09f14
          40725 => x"7f", -- $09f15
          40726 => x"7f", -- $09f16
          40727 => x"7f", -- $09f17
          40728 => x"7f", -- $09f18
          40729 => x"7f", -- $09f19
          40730 => x"7f", -- $09f1a
          40731 => x"7f", -- $09f1b
          40732 => x"7f", -- $09f1c
          40733 => x"7f", -- $09f1d
          40734 => x"7f", -- $09f1e
          40735 => x"7f", -- $09f1f
          40736 => x"7f", -- $09f20
          40737 => x"7f", -- $09f21
          40738 => x"7f", -- $09f22
          40739 => x"7f", -- $09f23
          40740 => x"7f", -- $09f24
          40741 => x"7f", -- $09f25
          40742 => x"7f", -- $09f26
          40743 => x"7f", -- $09f27
          40744 => x"7f", -- $09f28
          40745 => x"7f", -- $09f29
          40746 => x"7f", -- $09f2a
          40747 => x"7f", -- $09f2b
          40748 => x"7f", -- $09f2c
          40749 => x"7f", -- $09f2d
          40750 => x"7f", -- $09f2e
          40751 => x"7f", -- $09f2f
          40752 => x"7f", -- $09f30
          40753 => x"7f", -- $09f31
          40754 => x"7f", -- $09f32
          40755 => x"7f", -- $09f33
          40756 => x"7f", -- $09f34
          40757 => x"7f", -- $09f35
          40758 => x"7f", -- $09f36
          40759 => x"7f", -- $09f37
          40760 => x"7f", -- $09f38
          40761 => x"7f", -- $09f39
          40762 => x"7f", -- $09f3a
          40763 => x"7f", -- $09f3b
          40764 => x"7f", -- $09f3c
          40765 => x"7f", -- $09f3d
          40766 => x"7f", -- $09f3e
          40767 => x"7f", -- $09f3f
          40768 => x"7f", -- $09f40
          40769 => x"7f", -- $09f41
          40770 => x"7f", -- $09f42
          40771 => x"7f", -- $09f43
          40772 => x"7f", -- $09f44
          40773 => x"7f", -- $09f45
          40774 => x"7f", -- $09f46
          40775 => x"7f", -- $09f47
          40776 => x"7f", -- $09f48
          40777 => x"7f", -- $09f49
          40778 => x"7f", -- $09f4a
          40779 => x"7f", -- $09f4b
          40780 => x"7f", -- $09f4c
          40781 => x"7f", -- $09f4d
          40782 => x"7f", -- $09f4e
          40783 => x"7f", -- $09f4f
          40784 => x"7f", -- $09f50
          40785 => x"7f", -- $09f51
          40786 => x"7f", -- $09f52
          40787 => x"7f", -- $09f53
          40788 => x"7f", -- $09f54
          40789 => x"7f", -- $09f55
          40790 => x"7f", -- $09f56
          40791 => x"7f", -- $09f57
          40792 => x"7f", -- $09f58
          40793 => x"7f", -- $09f59
          40794 => x"7f", -- $09f5a
          40795 => x"7f", -- $09f5b
          40796 => x"7f", -- $09f5c
          40797 => x"7f", -- $09f5d
          40798 => x"7f", -- $09f5e
          40799 => x"7f", -- $09f5f
          40800 => x"7f", -- $09f60
          40801 => x"7f", -- $09f61
          40802 => x"7f", -- $09f62
          40803 => x"7f", -- $09f63
          40804 => x"7f", -- $09f64
          40805 => x"7f", -- $09f65
          40806 => x"7f", -- $09f66
          40807 => x"7f", -- $09f67
          40808 => x"7f", -- $09f68
          40809 => x"7f", -- $09f69
          40810 => x"7f", -- $09f6a
          40811 => x"7f", -- $09f6b
          40812 => x"7e", -- $09f6c
          40813 => x"7e", -- $09f6d
          40814 => x"7e", -- $09f6e
          40815 => x"7e", -- $09f6f
          40816 => x"7f", -- $09f70
          40817 => x"7f", -- $09f71
          40818 => x"7f", -- $09f72
          40819 => x"7f", -- $09f73
          40820 => x"7f", -- $09f74
          40821 => x"7e", -- $09f75
          40822 => x"7e", -- $09f76
          40823 => x"7e", -- $09f77
          40824 => x"7e", -- $09f78
          40825 => x"7e", -- $09f79
          40826 => x"7e", -- $09f7a
          40827 => x"7e", -- $09f7b
          40828 => x"7f", -- $09f7c
          40829 => x"7f", -- $09f7d
          40830 => x"7e", -- $09f7e
          40831 => x"7e", -- $09f7f
          40832 => x"7e", -- $09f80
          40833 => x"7e", -- $09f81
          40834 => x"7e", -- $09f82
          40835 => x"7e", -- $09f83
          40836 => x"7e", -- $09f84
          40837 => x"7e", -- $09f85
          40838 => x"7e", -- $09f86
          40839 => x"7e", -- $09f87
          40840 => x"7e", -- $09f88
          40841 => x"7e", -- $09f89
          40842 => x"7e", -- $09f8a
          40843 => x"7e", -- $09f8b
          40844 => x"7e", -- $09f8c
          40845 => x"7e", -- $09f8d
          40846 => x"7e", -- $09f8e
          40847 => x"7f", -- $09f8f
          40848 => x"7e", -- $09f90
          40849 => x"7e", -- $09f91
          40850 => x"7e", -- $09f92
          40851 => x"7e", -- $09f93
          40852 => x"7e", -- $09f94
          40853 => x"7e", -- $09f95
          40854 => x"7e", -- $09f96
          40855 => x"7e", -- $09f97
          40856 => x"7f", -- $09f98
          40857 => x"7f", -- $09f99
          40858 => x"7f", -- $09f9a
          40859 => x"7f", -- $09f9b
          40860 => x"7f", -- $09f9c
          40861 => x"7e", -- $09f9d
          40862 => x"7e", -- $09f9e
          40863 => x"7f", -- $09f9f
          40864 => x"7e", -- $09fa0
          40865 => x"7e", -- $09fa1
          40866 => x"7e", -- $09fa2
          40867 => x"7e", -- $09fa3
          40868 => x"7e", -- $09fa4
          40869 => x"7e", -- $09fa5
          40870 => x"7e", -- $09fa6
          40871 => x"7f", -- $09fa7
          40872 => x"7f", -- $09fa8
          40873 => x"7f", -- $09fa9
          40874 => x"7f", -- $09faa
          40875 => x"7f", -- $09fab
          40876 => x"7f", -- $09fac
          40877 => x"7f", -- $09fad
          40878 => x"7f", -- $09fae
          40879 => x"7f", -- $09faf
          40880 => x"7f", -- $09fb0
          40881 => x"7f", -- $09fb1
          40882 => x"7f", -- $09fb2
          40883 => x"7f", -- $09fb3
          40884 => x"7f", -- $09fb4
          40885 => x"7f", -- $09fb5
          40886 => x"7f", -- $09fb6
          40887 => x"7f", -- $09fb7
          40888 => x"7f", -- $09fb8
          40889 => x"7f", -- $09fb9
          40890 => x"7f", -- $09fba
          40891 => x"7f", -- $09fbb
          40892 => x"7f", -- $09fbc
          40893 => x"7f", -- $09fbd
          40894 => x"7f", -- $09fbe
          40895 => x"7f", -- $09fbf
          40896 => x"7f", -- $09fc0
          40897 => x"7f", -- $09fc1
          40898 => x"7f", -- $09fc2
          40899 => x"7f", -- $09fc3
          40900 => x"7f", -- $09fc4
          40901 => x"7f", -- $09fc5
          40902 => x"7f", -- $09fc6
          40903 => x"7f", -- $09fc7
          40904 => x"7f", -- $09fc8
          40905 => x"7f", -- $09fc9
          40906 => x"80", -- $09fca
          40907 => x"80", -- $09fcb
          40908 => x"80", -- $09fcc
          40909 => x"80", -- $09fcd
          40910 => x"80", -- $09fce
          40911 => x"80", -- $09fcf
          40912 => x"80", -- $09fd0
          40913 => x"80", -- $09fd1
          40914 => x"80", -- $09fd2
          40915 => x"80", -- $09fd3
          40916 => x"80", -- $09fd4
          40917 => x"80", -- $09fd5
          40918 => x"80", -- $09fd6
          40919 => x"7f", -- $09fd7
          40920 => x"7f", -- $09fd8
          40921 => x"7f", -- $09fd9
          40922 => x"7f", -- $09fda
          40923 => x"7f", -- $09fdb
          40924 => x"7f", -- $09fdc
          40925 => x"7f", -- $09fdd
          40926 => x"7f", -- $09fde
          40927 => x"80", -- $09fdf
          40928 => x"80", -- $09fe0
          40929 => x"80", -- $09fe1
          40930 => x"80", -- $09fe2
          40931 => x"80", -- $09fe3
          40932 => x"80", -- $09fe4
          40933 => x"80", -- $09fe5
          40934 => x"80", -- $09fe6
          40935 => x"80", -- $09fe7
          40936 => x"80", -- $09fe8
          40937 => x"80", -- $09fe9
          40938 => x"80", -- $09fea
          40939 => x"80", -- $09feb
          40940 => x"80", -- $09fec
          40941 => x"80", -- $09fed
          40942 => x"80", -- $09fee
          40943 => x"80", -- $09fef
          40944 => x"80", -- $09ff0
          40945 => x"80", -- $09ff1
          40946 => x"80", -- $09ff2
          40947 => x"80", -- $09ff3
          40948 => x"80", -- $09ff4
          40949 => x"80", -- $09ff5
          40950 => x"80", -- $09ff6
          40951 => x"80", -- $09ff7
          40952 => x"80", -- $09ff8
          40953 => x"80", -- $09ff9
          40954 => x"80", -- $09ffa
          40955 => x"80", -- $09ffb
          40956 => x"80", -- $09ffc
          40957 => x"80", -- $09ffd
          40958 => x"80", -- $09ffe
          40959 => x"80", -- $09fff
          40960 => x"80", -- $0a000
          40961 => x"80", -- $0a001
          40962 => x"80", -- $0a002
          40963 => x"80", -- $0a003
          40964 => x"80", -- $0a004
          40965 => x"80", -- $0a005
          40966 => x"80", -- $0a006
          40967 => x"80", -- $0a007
          40968 => x"80", -- $0a008
          40969 => x"80", -- $0a009
          40970 => x"80", -- $0a00a
          40971 => x"80", -- $0a00b
          40972 => x"80", -- $0a00c
          40973 => x"80", -- $0a00d
          40974 => x"80", -- $0a00e
          40975 => x"80", -- $0a00f
          40976 => x"80", -- $0a010
          40977 => x"80", -- $0a011
          40978 => x"80", -- $0a012
          40979 => x"80", -- $0a013
          40980 => x"80", -- $0a014
          40981 => x"80", -- $0a015
          40982 => x"80", -- $0a016
          40983 => x"80", -- $0a017
          40984 => x"80", -- $0a018
          40985 => x"80", -- $0a019
          40986 => x"80", -- $0a01a
          40987 => x"80", -- $0a01b
          40988 => x"80", -- $0a01c
          40989 => x"80", -- $0a01d
          40990 => x"80", -- $0a01e
          40991 => x"80", -- $0a01f
          40992 => x"80", -- $0a020
          40993 => x"80", -- $0a021
          40994 => x"80", -- $0a022
          40995 => x"80", -- $0a023
          40996 => x"80", -- $0a024
          40997 => x"80", -- $0a025
          40998 => x"80", -- $0a026
          40999 => x"80", -- $0a027
          41000 => x"80", -- $0a028
          41001 => x"80", -- $0a029
          41002 => x"80", -- $0a02a
          41003 => x"80", -- $0a02b
          41004 => x"80", -- $0a02c
          41005 => x"80", -- $0a02d
          41006 => x"80", -- $0a02e
          41007 => x"80", -- $0a02f
          41008 => x"80", -- $0a030
          41009 => x"80", -- $0a031
          41010 => x"80", -- $0a032
          41011 => x"80", -- $0a033
          41012 => x"80", -- $0a034
          41013 => x"81", -- $0a035
          41014 => x"81", -- $0a036
          41015 => x"81", -- $0a037
          41016 => x"81", -- $0a038
          41017 => x"81", -- $0a039
          41018 => x"81", -- $0a03a
          41019 => x"81", -- $0a03b
          41020 => x"81", -- $0a03c
          41021 => x"81", -- $0a03d
          41022 => x"81", -- $0a03e
          41023 => x"81", -- $0a03f
          41024 => x"80", -- $0a040
          41025 => x"80", -- $0a041
          41026 => x"80", -- $0a042
          41027 => x"80", -- $0a043
          41028 => x"80", -- $0a044
          41029 => x"80", -- $0a045
          41030 => x"80", -- $0a046
          41031 => x"80", -- $0a047
          41032 => x"80", -- $0a048
          41033 => x"80", -- $0a049
          41034 => x"80", -- $0a04a
          41035 => x"80", -- $0a04b
          41036 => x"80", -- $0a04c
          41037 => x"80", -- $0a04d
          41038 => x"81", -- $0a04e
          41039 => x"81", -- $0a04f
          41040 => x"81", -- $0a050
          41041 => x"81", -- $0a051
          41042 => x"81", -- $0a052
          41043 => x"81", -- $0a053
          41044 => x"81", -- $0a054
          41045 => x"81", -- $0a055
          41046 => x"81", -- $0a056
          41047 => x"81", -- $0a057
          41048 => x"81", -- $0a058
          41049 => x"81", -- $0a059
          41050 => x"81", -- $0a05a
          41051 => x"81", -- $0a05b
          41052 => x"81", -- $0a05c
          41053 => x"81", -- $0a05d
          41054 => x"80", -- $0a05e
          41055 => x"80", -- $0a05f
          41056 => x"80", -- $0a060
          41057 => x"80", -- $0a061
          41058 => x"80", -- $0a062
          41059 => x"80", -- $0a063
          41060 => x"80", -- $0a064
          41061 => x"81", -- $0a065
          41062 => x"81", -- $0a066
          41063 => x"81", -- $0a067
          41064 => x"81", -- $0a068
          41065 => x"81", -- $0a069
          41066 => x"81", -- $0a06a
          41067 => x"81", -- $0a06b
          41068 => x"81", -- $0a06c
          41069 => x"81", -- $0a06d
          41070 => x"81", -- $0a06e
          41071 => x"81", -- $0a06f
          41072 => x"81", -- $0a070
          41073 => x"81", -- $0a071
          41074 => x"81", -- $0a072
          41075 => x"81", -- $0a073
          41076 => x"81", -- $0a074
          41077 => x"81", -- $0a075
          41078 => x"81", -- $0a076
          41079 => x"81", -- $0a077
          41080 => x"81", -- $0a078
          41081 => x"81", -- $0a079
          41082 => x"81", -- $0a07a
          41083 => x"81", -- $0a07b
          41084 => x"81", -- $0a07c
          41085 => x"81", -- $0a07d
          41086 => x"81", -- $0a07e
          41087 => x"81", -- $0a07f
          41088 => x"81", -- $0a080
          41089 => x"81", -- $0a081
          41090 => x"81", -- $0a082
          41091 => x"81", -- $0a083
          41092 => x"81", -- $0a084
          41093 => x"81", -- $0a085
          41094 => x"82", -- $0a086
          41095 => x"81", -- $0a087
          41096 => x"81", -- $0a088
          41097 => x"81", -- $0a089
          41098 => x"81", -- $0a08a
          41099 => x"81", -- $0a08b
          41100 => x"81", -- $0a08c
          41101 => x"81", -- $0a08d
          41102 => x"81", -- $0a08e
          41103 => x"81", -- $0a08f
          41104 => x"81", -- $0a090
          41105 => x"81", -- $0a091
          41106 => x"81", -- $0a092
          41107 => x"81", -- $0a093
          41108 => x"81", -- $0a094
          41109 => x"80", -- $0a095
          41110 => x"81", -- $0a096
          41111 => x"81", -- $0a097
          41112 => x"81", -- $0a098
          41113 => x"81", -- $0a099
          41114 => x"81", -- $0a09a
          41115 => x"81", -- $0a09b
          41116 => x"81", -- $0a09c
          41117 => x"81", -- $0a09d
          41118 => x"81", -- $0a09e
          41119 => x"81", -- $0a09f
          41120 => x"82", -- $0a0a0
          41121 => x"81", -- $0a0a1
          41122 => x"81", -- $0a0a2
          41123 => x"81", -- $0a0a3
          41124 => x"81", -- $0a0a4
          41125 => x"81", -- $0a0a5
          41126 => x"81", -- $0a0a6
          41127 => x"81", -- $0a0a7
          41128 => x"81", -- $0a0a8
          41129 => x"81", -- $0a0a9
          41130 => x"81", -- $0a0aa
          41131 => x"81", -- $0a0ab
          41132 => x"81", -- $0a0ac
          41133 => x"81", -- $0a0ad
          41134 => x"81", -- $0a0ae
          41135 => x"81", -- $0a0af
          41136 => x"81", -- $0a0b0
          41137 => x"81", -- $0a0b1
          41138 => x"81", -- $0a0b2
          41139 => x"81", -- $0a0b3
          41140 => x"81", -- $0a0b4
          41141 => x"81", -- $0a0b5
          41142 => x"81", -- $0a0b6
          41143 => x"82", -- $0a0b7
          41144 => x"82", -- $0a0b8
          41145 => x"82", -- $0a0b9
          41146 => x"82", -- $0a0ba
          41147 => x"82", -- $0a0bb
          41148 => x"82", -- $0a0bc
          41149 => x"82", -- $0a0bd
          41150 => x"82", -- $0a0be
          41151 => x"82", -- $0a0bf
          41152 => x"81", -- $0a0c0
          41153 => x"81", -- $0a0c1
          41154 => x"81", -- $0a0c2
          41155 => x"81", -- $0a0c3
          41156 => x"81", -- $0a0c4
          41157 => x"81", -- $0a0c5
          41158 => x"81", -- $0a0c6
          41159 => x"81", -- $0a0c7
          41160 => x"81", -- $0a0c8
          41161 => x"81", -- $0a0c9
          41162 => x"81", -- $0a0ca
          41163 => x"81", -- $0a0cb
          41164 => x"81", -- $0a0cc
          41165 => x"81", -- $0a0cd
          41166 => x"82", -- $0a0ce
          41167 => x"82", -- $0a0cf
          41168 => x"82", -- $0a0d0
          41169 => x"82", -- $0a0d1
          41170 => x"82", -- $0a0d2
          41171 => x"82", -- $0a0d3
          41172 => x"82", -- $0a0d4
          41173 => x"82", -- $0a0d5
          41174 => x"82", -- $0a0d6
          41175 => x"82", -- $0a0d7
          41176 => x"82", -- $0a0d8
          41177 => x"82", -- $0a0d9
          41178 => x"82", -- $0a0da
          41179 => x"82", -- $0a0db
          41180 => x"82", -- $0a0dc
          41181 => x"81", -- $0a0dd
          41182 => x"81", -- $0a0de
          41183 => x"81", -- $0a0df
          41184 => x"81", -- $0a0e0
          41185 => x"81", -- $0a0e1
          41186 => x"81", -- $0a0e2
          41187 => x"81", -- $0a0e3
          41188 => x"81", -- $0a0e4
          41189 => x"81", -- $0a0e5
          41190 => x"81", -- $0a0e6
          41191 => x"82", -- $0a0e7
          41192 => x"82", -- $0a0e8
          41193 => x"82", -- $0a0e9
          41194 => x"82", -- $0a0ea
          41195 => x"82", -- $0a0eb
          41196 => x"82", -- $0a0ec
          41197 => x"82", -- $0a0ed
          41198 => x"82", -- $0a0ee
          41199 => x"82", -- $0a0ef
          41200 => x"82", -- $0a0f0
          41201 => x"82", -- $0a0f1
          41202 => x"82", -- $0a0f2
          41203 => x"82", -- $0a0f3
          41204 => x"82", -- $0a0f4
          41205 => x"82", -- $0a0f5
          41206 => x"82", -- $0a0f6
          41207 => x"81", -- $0a0f7
          41208 => x"81", -- $0a0f8
          41209 => x"81", -- $0a0f9
          41210 => x"81", -- $0a0fa
          41211 => x"81", -- $0a0fb
          41212 => x"81", -- $0a0fc
          41213 => x"81", -- $0a0fd
          41214 => x"81", -- $0a0fe
          41215 => x"81", -- $0a0ff
          41216 => x"81", -- $0a100
          41217 => x"81", -- $0a101
          41218 => x"81", -- $0a102
          41219 => x"82", -- $0a103
          41220 => x"82", -- $0a104
          41221 => x"82", -- $0a105
          41222 => x"82", -- $0a106
          41223 => x"82", -- $0a107
          41224 => x"82", -- $0a108
          41225 => x"82", -- $0a109
          41226 => x"82", -- $0a10a
          41227 => x"82", -- $0a10b
          41228 => x"82", -- $0a10c
          41229 => x"82", -- $0a10d
          41230 => x"82", -- $0a10e
          41231 => x"81", -- $0a10f
          41232 => x"81", -- $0a110
          41233 => x"81", -- $0a111
          41234 => x"81", -- $0a112
          41235 => x"81", -- $0a113
          41236 => x"80", -- $0a114
          41237 => x"80", -- $0a115
          41238 => x"80", -- $0a116
          41239 => x"80", -- $0a117
          41240 => x"80", -- $0a118
          41241 => x"81", -- $0a119
          41242 => x"81", -- $0a11a
          41243 => x"81", -- $0a11b
          41244 => x"81", -- $0a11c
          41245 => x"81", -- $0a11d
          41246 => x"81", -- $0a11e
          41247 => x"81", -- $0a11f
          41248 => x"81", -- $0a120
          41249 => x"82", -- $0a121
          41250 => x"82", -- $0a122
          41251 => x"82", -- $0a123
          41252 => x"82", -- $0a124
          41253 => x"82", -- $0a125
          41254 => x"82", -- $0a126
          41255 => x"81", -- $0a127
          41256 => x"81", -- $0a128
          41257 => x"81", -- $0a129
          41258 => x"81", -- $0a12a
          41259 => x"80", -- $0a12b
          41260 => x"80", -- $0a12c
          41261 => x"80", -- $0a12d
          41262 => x"80", -- $0a12e
          41263 => x"80", -- $0a12f
          41264 => x"80", -- $0a130
          41265 => x"80", -- $0a131
          41266 => x"80", -- $0a132
          41267 => x"80", -- $0a133
          41268 => x"80", -- $0a134
          41269 => x"80", -- $0a135
          41270 => x"80", -- $0a136
          41271 => x"80", -- $0a137
          41272 => x"80", -- $0a138
          41273 => x"81", -- $0a139
          41274 => x"81", -- $0a13a
          41275 => x"81", -- $0a13b
          41276 => x"81", -- $0a13c
          41277 => x"81", -- $0a13d
          41278 => x"81", -- $0a13e
          41279 => x"81", -- $0a13f
          41280 => x"81", -- $0a140
          41281 => x"81", -- $0a141
          41282 => x"81", -- $0a142
          41283 => x"80", -- $0a143
          41284 => x"80", -- $0a144
          41285 => x"80", -- $0a145
          41286 => x"80", -- $0a146
          41287 => x"80", -- $0a147
          41288 => x"80", -- $0a148
          41289 => x"80", -- $0a149
          41290 => x"80", -- $0a14a
          41291 => x"80", -- $0a14b
          41292 => x"80", -- $0a14c
          41293 => x"80", -- $0a14d
          41294 => x"80", -- $0a14e
          41295 => x"80", -- $0a14f
          41296 => x"80", -- $0a150
          41297 => x"80", -- $0a151
          41298 => x"80", -- $0a152
          41299 => x"80", -- $0a153
          41300 => x"80", -- $0a154
          41301 => x"80", -- $0a155
          41302 => x"80", -- $0a156
          41303 => x"80", -- $0a157
          41304 => x"81", -- $0a158
          41305 => x"80", -- $0a159
          41306 => x"80", -- $0a15a
          41307 => x"80", -- $0a15b
          41308 => x"80", -- $0a15c
          41309 => x"80", -- $0a15d
          41310 => x"80", -- $0a15e
          41311 => x"80", -- $0a15f
          41312 => x"80", -- $0a160
          41313 => x"80", -- $0a161
          41314 => x"80", -- $0a162
          41315 => x"80", -- $0a163
          41316 => x"80", -- $0a164
          41317 => x"80", -- $0a165
          41318 => x"80", -- $0a166
          41319 => x"80", -- $0a167
          41320 => x"80", -- $0a168
          41321 => x"80", -- $0a169
          41322 => x"80", -- $0a16a
          41323 => x"80", -- $0a16b
          41324 => x"80", -- $0a16c
          41325 => x"80", -- $0a16d
          41326 => x"80", -- $0a16e
          41327 => x"80", -- $0a16f
          41328 => x"80", -- $0a170
          41329 => x"80", -- $0a171
          41330 => x"80", -- $0a172
          41331 => x"80", -- $0a173
          41332 => x"80", -- $0a174
          41333 => x"80", -- $0a175
          41334 => x"80", -- $0a176
          41335 => x"80", -- $0a177
          41336 => x"80", -- $0a178
          41337 => x"80", -- $0a179
          41338 => x"80", -- $0a17a
          41339 => x"80", -- $0a17b
          41340 => x"7f", -- $0a17c
          41341 => x"7f", -- $0a17d
          41342 => x"7f", -- $0a17e
          41343 => x"7f", -- $0a17f
          41344 => x"7f", -- $0a180
          41345 => x"7f", -- $0a181
          41346 => x"7f", -- $0a182
          41347 => x"7f", -- $0a183
          41348 => x"7f", -- $0a184
          41349 => x"80", -- $0a185
          41350 => x"80", -- $0a186
          41351 => x"80", -- $0a187
          41352 => x"80", -- $0a188
          41353 => x"80", -- $0a189
          41354 => x"80", -- $0a18a
          41355 => x"80", -- $0a18b
          41356 => x"80", -- $0a18c
          41357 => x"80", -- $0a18d
          41358 => x"80", -- $0a18e
          41359 => x"80", -- $0a18f
          41360 => x"80", -- $0a190
          41361 => x"80", -- $0a191
          41362 => x"80", -- $0a192
          41363 => x"7f", -- $0a193
          41364 => x"7f", -- $0a194
          41365 => x"7f", -- $0a195
          41366 => x"7f", -- $0a196
          41367 => x"7f", -- $0a197
          41368 => x"7f", -- $0a198
          41369 => x"7f", -- $0a199
          41370 => x"7f", -- $0a19a
          41371 => x"7f", -- $0a19b
          41372 => x"7f", -- $0a19c
          41373 => x"7f", -- $0a19d
          41374 => x"7f", -- $0a19e
          41375 => x"7f", -- $0a19f
          41376 => x"80", -- $0a1a0
          41377 => x"80", -- $0a1a1
          41378 => x"80", -- $0a1a2
          41379 => x"80", -- $0a1a3
          41380 => x"80", -- $0a1a4
          41381 => x"80", -- $0a1a5
          41382 => x"80", -- $0a1a6
          41383 => x"80", -- $0a1a7
          41384 => x"80", -- $0a1a8
          41385 => x"80", -- $0a1a9
          41386 => x"80", -- $0a1aa
          41387 => x"80", -- $0a1ab
          41388 => x"7f", -- $0a1ac
          41389 => x"7f", -- $0a1ad
          41390 => x"7f", -- $0a1ae
          41391 => x"7f", -- $0a1af
          41392 => x"7f", -- $0a1b0
          41393 => x"7f", -- $0a1b1
          41394 => x"7f", -- $0a1b2
          41395 => x"7f", -- $0a1b3
          41396 => x"7f", -- $0a1b4
          41397 => x"7f", -- $0a1b5
          41398 => x"7f", -- $0a1b6
          41399 => x"7f", -- $0a1b7
          41400 => x"7f", -- $0a1b8
          41401 => x"7f", -- $0a1b9
          41402 => x"7f", -- $0a1ba
          41403 => x"80", -- $0a1bb
          41404 => x"80", -- $0a1bc
          41405 => x"80", -- $0a1bd
          41406 => x"80", -- $0a1be
          41407 => x"80", -- $0a1bf
          41408 => x"80", -- $0a1c0
          41409 => x"80", -- $0a1c1
          41410 => x"80", -- $0a1c2
          41411 => x"80", -- $0a1c3
          41412 => x"80", -- $0a1c4
          41413 => x"7f", -- $0a1c5
          41414 => x"7f", -- $0a1c6
          41415 => x"7f", -- $0a1c7
          41416 => x"7f", -- $0a1c8
          41417 => x"7f", -- $0a1c9
          41418 => x"7f", -- $0a1ca
          41419 => x"7f", -- $0a1cb
          41420 => x"7f", -- $0a1cc
          41421 => x"7f", -- $0a1cd
          41422 => x"7f", -- $0a1ce
          41423 => x"7f", -- $0a1cf
          41424 => x"7f", -- $0a1d0
          41425 => x"7f", -- $0a1d1
          41426 => x"7f", -- $0a1d2
          41427 => x"7f", -- $0a1d3
          41428 => x"7f", -- $0a1d4
          41429 => x"7f", -- $0a1d5
          41430 => x"80", -- $0a1d6
          41431 => x"80", -- $0a1d7
          41432 => x"80", -- $0a1d8
          41433 => x"80", -- $0a1d9
          41434 => x"80", -- $0a1da
          41435 => x"80", -- $0a1db
          41436 => x"80", -- $0a1dc
          41437 => x"7f", -- $0a1dd
          41438 => x"7f", -- $0a1de
          41439 => x"7f", -- $0a1df
          41440 => x"7f", -- $0a1e0
          41441 => x"7e", -- $0a1e1
          41442 => x"7e", -- $0a1e2
          41443 => x"7e", -- $0a1e3
          41444 => x"7e", -- $0a1e4
          41445 => x"7e", -- $0a1e5
          41446 => x"7e", -- $0a1e6
          41447 => x"7e", -- $0a1e7
          41448 => x"7e", -- $0a1e8
          41449 => x"7e", -- $0a1e9
          41450 => x"7e", -- $0a1ea
          41451 => x"7e", -- $0a1eb
          41452 => x"7e", -- $0a1ec
          41453 => x"7f", -- $0a1ed
          41454 => x"7f", -- $0a1ee
          41455 => x"7f", -- $0a1ef
          41456 => x"7f", -- $0a1f0
          41457 => x"7f", -- $0a1f1
          41458 => x"7f", -- $0a1f2
          41459 => x"7f", -- $0a1f3
          41460 => x"7f", -- $0a1f4
          41461 => x"7f", -- $0a1f5
          41462 => x"7f", -- $0a1f6
          41463 => x"7f", -- $0a1f7
          41464 => x"7f", -- $0a1f8
          41465 => x"7f", -- $0a1f9
          41466 => x"7f", -- $0a1fa
          41467 => x"7e", -- $0a1fb
          41468 => x"7e", -- $0a1fc
          41469 => x"7e", -- $0a1fd
          41470 => x"7e", -- $0a1fe
          41471 => x"7e", -- $0a1ff
          41472 => x"7e", -- $0a200
          41473 => x"7e", -- $0a201
          41474 => x"7e", -- $0a202
          41475 => x"7e", -- $0a203
          41476 => x"7e", -- $0a204
          41477 => x"7e", -- $0a205
          41478 => x"7e", -- $0a206
          41479 => x"7e", -- $0a207
          41480 => x"7e", -- $0a208
          41481 => x"7f", -- $0a209
          41482 => x"7f", -- $0a20a
          41483 => x"7f", -- $0a20b
          41484 => x"7f", -- $0a20c
          41485 => x"7f", -- $0a20d
          41486 => x"7f", -- $0a20e
          41487 => x"7f", -- $0a20f
          41488 => x"7f", -- $0a210
          41489 => x"7f", -- $0a211
          41490 => x"7f", -- $0a212
          41491 => x"7f", -- $0a213
          41492 => x"7e", -- $0a214
          41493 => x"7e", -- $0a215
          41494 => x"7e", -- $0a216
          41495 => x"7e", -- $0a217
          41496 => x"7e", -- $0a218
          41497 => x"7e", -- $0a219
          41498 => x"7e", -- $0a21a
          41499 => x"7e", -- $0a21b
          41500 => x"7e", -- $0a21c
          41501 => x"7e", -- $0a21d
          41502 => x"7e", -- $0a21e
          41503 => x"7e", -- $0a21f
          41504 => x"7e", -- $0a220
          41505 => x"7e", -- $0a221
          41506 => x"7e", -- $0a222
          41507 => x"7f", -- $0a223
          41508 => x"7f", -- $0a224
          41509 => x"7f", -- $0a225
          41510 => x"7f", -- $0a226
          41511 => x"7f", -- $0a227
          41512 => x"7f", -- $0a228
          41513 => x"7f", -- $0a229
          41514 => x"7f", -- $0a22a
          41515 => x"7f", -- $0a22b
          41516 => x"7f", -- $0a22c
          41517 => x"7f", -- $0a22d
          41518 => x"7f", -- $0a22e
          41519 => x"7f", -- $0a22f
          41520 => x"7f", -- $0a230
          41521 => x"7f", -- $0a231
          41522 => x"7f", -- $0a232
          41523 => x"7e", -- $0a233
          41524 => x"7e", -- $0a234
          41525 => x"7e", -- $0a235
          41526 => x"7e", -- $0a236
          41527 => x"7e", -- $0a237
          41528 => x"7e", -- $0a238
          41529 => x"7e", -- $0a239
          41530 => x"7e", -- $0a23a
          41531 => x"7e", -- $0a23b
          41532 => x"7f", -- $0a23c
          41533 => x"7f", -- $0a23d
          41534 => x"7f", -- $0a23e
          41535 => x"7f", -- $0a23f
          41536 => x"7f", -- $0a240
          41537 => x"7f", -- $0a241
          41538 => x"7f", -- $0a242
          41539 => x"7f", -- $0a243
          41540 => x"7f", -- $0a244
          41541 => x"7f", -- $0a245
          41542 => x"7f", -- $0a246
          41543 => x"7f", -- $0a247
          41544 => x"7f", -- $0a248
          41545 => x"7f", -- $0a249
          41546 => x"7f", -- $0a24a
          41547 => x"7f", -- $0a24b
          41548 => x"7f", -- $0a24c
          41549 => x"7f", -- $0a24d
          41550 => x"7e", -- $0a24e
          41551 => x"7e", -- $0a24f
          41552 => x"7e", -- $0a250
          41553 => x"7e", -- $0a251
          41554 => x"7e", -- $0a252
          41555 => x"7e", -- $0a253
          41556 => x"7e", -- $0a254
          41557 => x"7e", -- $0a255
          41558 => x"7e", -- $0a256
          41559 => x"7f", -- $0a257
          41560 => x"7f", -- $0a258
          41561 => x"7f", -- $0a259
          41562 => x"7f", -- $0a25a
          41563 => x"7f", -- $0a25b
          41564 => x"7f", -- $0a25c
          41565 => x"7f", -- $0a25d
          41566 => x"7f", -- $0a25e
          41567 => x"7f", -- $0a25f
          41568 => x"7f", -- $0a260
          41569 => x"7f", -- $0a261
          41570 => x"7f", -- $0a262
          41571 => x"7f", -- $0a263
          41572 => x"7f", -- $0a264
          41573 => x"7f", -- $0a265
          41574 => x"7f", -- $0a266
          41575 => x"7f", -- $0a267
          41576 => x"7f", -- $0a268
          41577 => x"7f", -- $0a269
          41578 => x"7e", -- $0a26a
          41579 => x"7e", -- $0a26b
          41580 => x"7e", -- $0a26c
          41581 => x"7e", -- $0a26d
          41582 => x"7f", -- $0a26e
          41583 => x"7f", -- $0a26f
          41584 => x"7f", -- $0a270
          41585 => x"7f", -- $0a271
          41586 => x"7f", -- $0a272
          41587 => x"7f", -- $0a273
          41588 => x"7f", -- $0a274
          41589 => x"7f", -- $0a275
          41590 => x"7f", -- $0a276
          41591 => x"7f", -- $0a277
          41592 => x"7f", -- $0a278
          41593 => x"7f", -- $0a279
          41594 => x"7f", -- $0a27a
          41595 => x"7f", -- $0a27b
          41596 => x"7f", -- $0a27c
          41597 => x"7f", -- $0a27d
          41598 => x"7f", -- $0a27e
          41599 => x"7f", -- $0a27f
          41600 => x"7f", -- $0a280
          41601 => x"7f", -- $0a281
          41602 => x"7f", -- $0a282
          41603 => x"7f", -- $0a283
          41604 => x"7f", -- $0a284
          41605 => x"7f", -- $0a285
          41606 => x"7f", -- $0a286
          41607 => x"7f", -- $0a287
          41608 => x"7f", -- $0a288
          41609 => x"7f", -- $0a289
          41610 => x"7f", -- $0a28a
          41611 => x"7f", -- $0a28b
          41612 => x"7f", -- $0a28c
          41613 => x"7f", -- $0a28d
          41614 => x"7f", -- $0a28e
          41615 => x"80", -- $0a28f
          41616 => x"80", -- $0a290
          41617 => x"80", -- $0a291
          41618 => x"80", -- $0a292
          41619 => x"7f", -- $0a293
          41620 => x"7f", -- $0a294
          41621 => x"7f", -- $0a295
          41622 => x"80", -- $0a296
          41623 => x"7f", -- $0a297
          41624 => x"7f", -- $0a298
          41625 => x"7f", -- $0a299
          41626 => x"7f", -- $0a29a
          41627 => x"7f", -- $0a29b
          41628 => x"7f", -- $0a29c
          41629 => x"7f", -- $0a29d
          41630 => x"7f", -- $0a29e
          41631 => x"7f", -- $0a29f
          41632 => x"7f", -- $0a2a0
          41633 => x"7f", -- $0a2a1
          41634 => x"7f", -- $0a2a2
          41635 => x"7f", -- $0a2a3
          41636 => x"7f", -- $0a2a4
          41637 => x"80", -- $0a2a5
          41638 => x"80", -- $0a2a6
          41639 => x"80", -- $0a2a7
          41640 => x"80", -- $0a2a8
          41641 => x"80", -- $0a2a9
          41642 => x"80", -- $0a2aa
          41643 => x"80", -- $0a2ab
          41644 => x"80", -- $0a2ac
          41645 => x"80", -- $0a2ad
          41646 => x"80", -- $0a2ae
          41647 => x"80", -- $0a2af
          41648 => x"7f", -- $0a2b0
          41649 => x"80", -- $0a2b1
          41650 => x"80", -- $0a2b2
          41651 => x"7f", -- $0a2b3
          41652 => x"7f", -- $0a2b4
          41653 => x"7f", -- $0a2b5
          41654 => x"7f", -- $0a2b6
          41655 => x"7f", -- $0a2b7
          41656 => x"7f", -- $0a2b8
          41657 => x"7f", -- $0a2b9
          41658 => x"80", -- $0a2ba
          41659 => x"80", -- $0a2bb
          41660 => x"80", -- $0a2bc
          41661 => x"80", -- $0a2bd
          41662 => x"80", -- $0a2be
          41663 => x"80", -- $0a2bf
          41664 => x"80", -- $0a2c0
          41665 => x"80", -- $0a2c1
          41666 => x"80", -- $0a2c2
          41667 => x"80", -- $0a2c3
          41668 => x"80", -- $0a2c4
          41669 => x"80", -- $0a2c5
          41670 => x"80", -- $0a2c6
          41671 => x"80", -- $0a2c7
          41672 => x"80", -- $0a2c8
          41673 => x"80", -- $0a2c9
          41674 => x"80", -- $0a2ca
          41675 => x"80", -- $0a2cb
          41676 => x"80", -- $0a2cc
          41677 => x"80", -- $0a2cd
          41678 => x"80", -- $0a2ce
          41679 => x"80", -- $0a2cf
          41680 => x"80", -- $0a2d0
          41681 => x"80", -- $0a2d1
          41682 => x"80", -- $0a2d2
          41683 => x"80", -- $0a2d3
          41684 => x"80", -- $0a2d4
          41685 => x"80", -- $0a2d5
          41686 => x"80", -- $0a2d6
          41687 => x"80", -- $0a2d7
          41688 => x"80", -- $0a2d8
          41689 => x"80", -- $0a2d9
          41690 => x"80", -- $0a2da
          41691 => x"80", -- $0a2db
          41692 => x"80", -- $0a2dc
          41693 => x"80", -- $0a2dd
          41694 => x"80", -- $0a2de
          41695 => x"80", -- $0a2df
          41696 => x"80", -- $0a2e0
          41697 => x"80", -- $0a2e1
          41698 => x"80", -- $0a2e2
          41699 => x"80", -- $0a2e3
          41700 => x"80", -- $0a2e4
          41701 => x"80", -- $0a2e5
          41702 => x"80", -- $0a2e6
          41703 => x"80", -- $0a2e7
          41704 => x"80", -- $0a2e8
          41705 => x"80", -- $0a2e9
          41706 => x"80", -- $0a2ea
          41707 => x"80", -- $0a2eb
          41708 => x"80", -- $0a2ec
          41709 => x"80", -- $0a2ed
          41710 => x"80", -- $0a2ee
          41711 => x"80", -- $0a2ef
          41712 => x"80", -- $0a2f0
          41713 => x"80", -- $0a2f1
          41714 => x"80", -- $0a2f2
          41715 => x"80", -- $0a2f3
          41716 => x"80", -- $0a2f4
          41717 => x"80", -- $0a2f5
          41718 => x"80", -- $0a2f6
          41719 => x"80", -- $0a2f7
          41720 => x"80", -- $0a2f8
          41721 => x"80", -- $0a2f9
          41722 => x"80", -- $0a2fa
          41723 => x"80", -- $0a2fb
          41724 => x"80", -- $0a2fc
          41725 => x"80", -- $0a2fd
          41726 => x"80", -- $0a2fe
          41727 => x"80", -- $0a2ff
          41728 => x"80", -- $0a300
          41729 => x"80", -- $0a301
          41730 => x"80", -- $0a302
          41731 => x"80", -- $0a303
          41732 => x"80", -- $0a304
          41733 => x"80", -- $0a305
          41734 => x"80", -- $0a306
          41735 => x"80", -- $0a307
          41736 => x"80", -- $0a308
          41737 => x"80", -- $0a309
          41738 => x"80", -- $0a30a
          41739 => x"80", -- $0a30b
          41740 => x"80", -- $0a30c
          41741 => x"80", -- $0a30d
          41742 => x"80", -- $0a30e
          41743 => x"81", -- $0a30f
          41744 => x"81", -- $0a310
          41745 => x"81", -- $0a311
          41746 => x"81", -- $0a312
          41747 => x"81", -- $0a313
          41748 => x"81", -- $0a314
          41749 => x"80", -- $0a315
          41750 => x"80", -- $0a316
          41751 => x"80", -- $0a317
          41752 => x"80", -- $0a318
          41753 => x"80", -- $0a319
          41754 => x"80", -- $0a31a
          41755 => x"80", -- $0a31b
          41756 => x"80", -- $0a31c
          41757 => x"80", -- $0a31d
          41758 => x"80", -- $0a31e
          41759 => x"80", -- $0a31f
          41760 => x"80", -- $0a320
          41761 => x"80", -- $0a321
          41762 => x"80", -- $0a322
          41763 => x"80", -- $0a323
          41764 => x"80", -- $0a324
          41765 => x"80", -- $0a325
          41766 => x"80", -- $0a326
          41767 => x"81", -- $0a327
          41768 => x"81", -- $0a328
          41769 => x"81", -- $0a329
          41770 => x"81", -- $0a32a
          41771 => x"81", -- $0a32b
          41772 => x"81", -- $0a32c
          41773 => x"81", -- $0a32d
          41774 => x"81", -- $0a32e
          41775 => x"81", -- $0a32f
          41776 => x"81", -- $0a330
          41777 => x"81", -- $0a331
          41778 => x"81", -- $0a332
          41779 => x"81", -- $0a333
          41780 => x"81", -- $0a334
          41781 => x"81", -- $0a335
          41782 => x"81", -- $0a336
          41783 => x"81", -- $0a337
          41784 => x"81", -- $0a338
          41785 => x"81", -- $0a339
          41786 => x"81", -- $0a33a
          41787 => x"81", -- $0a33b
          41788 => x"81", -- $0a33c
          41789 => x"81", -- $0a33d
          41790 => x"81", -- $0a33e
          41791 => x"81", -- $0a33f
          41792 => x"81", -- $0a340
          41793 => x"81", -- $0a341
          41794 => x"81", -- $0a342
          41795 => x"81", -- $0a343
          41796 => x"81", -- $0a344
          41797 => x"81", -- $0a345
          41798 => x"81", -- $0a346
          41799 => x"81", -- $0a347
          41800 => x"81", -- $0a348
          41801 => x"81", -- $0a349
          41802 => x"81", -- $0a34a
          41803 => x"81", -- $0a34b
          41804 => x"81", -- $0a34c
          41805 => x"81", -- $0a34d
          41806 => x"81", -- $0a34e
          41807 => x"81", -- $0a34f
          41808 => x"81", -- $0a350
          41809 => x"81", -- $0a351
          41810 => x"81", -- $0a352
          41811 => x"81", -- $0a353
          41812 => x"81", -- $0a354
          41813 => x"81", -- $0a355
          41814 => x"81", -- $0a356
          41815 => x"81", -- $0a357
          41816 => x"81", -- $0a358
          41817 => x"81", -- $0a359
          41818 => x"82", -- $0a35a
          41819 => x"82", -- $0a35b
          41820 => x"82", -- $0a35c
          41821 => x"82", -- $0a35d
          41822 => x"82", -- $0a35e
          41823 => x"82", -- $0a35f
          41824 => x"82", -- $0a360
          41825 => x"82", -- $0a361
          41826 => x"82", -- $0a362
          41827 => x"82", -- $0a363
          41828 => x"82", -- $0a364
          41829 => x"82", -- $0a365
          41830 => x"82", -- $0a366
          41831 => x"82", -- $0a367
          41832 => x"82", -- $0a368
          41833 => x"82", -- $0a369
          41834 => x"82", -- $0a36a
          41835 => x"82", -- $0a36b
          41836 => x"81", -- $0a36c
          41837 => x"82", -- $0a36d
          41838 => x"82", -- $0a36e
          41839 => x"81", -- $0a36f
          41840 => x"82", -- $0a370
          41841 => x"82", -- $0a371
          41842 => x"82", -- $0a372
          41843 => x"82", -- $0a373
          41844 => x"82", -- $0a374
          41845 => x"82", -- $0a375
          41846 => x"82", -- $0a376
          41847 => x"82", -- $0a377
          41848 => x"82", -- $0a378
          41849 => x"82", -- $0a379
          41850 => x"82", -- $0a37a
          41851 => x"82", -- $0a37b
          41852 => x"82", -- $0a37c
          41853 => x"82", -- $0a37d
          41854 => x"82", -- $0a37e
          41855 => x"82", -- $0a37f
          41856 => x"82", -- $0a380
          41857 => x"82", -- $0a381
          41858 => x"82", -- $0a382
          41859 => x"82", -- $0a383
          41860 => x"82", -- $0a384
          41861 => x"82", -- $0a385
          41862 => x"82", -- $0a386
          41863 => x"82", -- $0a387
          41864 => x"82", -- $0a388
          41865 => x"82", -- $0a389
          41866 => x"82", -- $0a38a
          41867 => x"82", -- $0a38b
          41868 => x"82", -- $0a38c
          41869 => x"82", -- $0a38d
          41870 => x"82", -- $0a38e
          41871 => x"82", -- $0a38f
          41872 => x"82", -- $0a390
          41873 => x"82", -- $0a391
          41874 => x"82", -- $0a392
          41875 => x"82", -- $0a393
          41876 => x"82", -- $0a394
          41877 => x"82", -- $0a395
          41878 => x"82", -- $0a396
          41879 => x"82", -- $0a397
          41880 => x"82", -- $0a398
          41881 => x"82", -- $0a399
          41882 => x"82", -- $0a39a
          41883 => x"81", -- $0a39b
          41884 => x"81", -- $0a39c
          41885 => x"81", -- $0a39d
          41886 => x"81", -- $0a39e
          41887 => x"81", -- $0a39f
          41888 => x"81", -- $0a3a0
          41889 => x"81", -- $0a3a1
          41890 => x"81", -- $0a3a2
          41891 => x"81", -- $0a3a3
          41892 => x"81", -- $0a3a4
          41893 => x"81", -- $0a3a5
          41894 => x"81", -- $0a3a6
          41895 => x"81", -- $0a3a7
          41896 => x"81", -- $0a3a8
          41897 => x"81", -- $0a3a9
          41898 => x"81", -- $0a3aa
          41899 => x"81", -- $0a3ab
          41900 => x"81", -- $0a3ac
          41901 => x"81", -- $0a3ad
          41902 => x"81", -- $0a3ae
          41903 => x"81", -- $0a3af
          41904 => x"81", -- $0a3b0
          41905 => x"81", -- $0a3b1
          41906 => x"81", -- $0a3b2
          41907 => x"81", -- $0a3b3
          41908 => x"81", -- $0a3b4
          41909 => x"81", -- $0a3b5
          41910 => x"81", -- $0a3b6
          41911 => x"81", -- $0a3b7
          41912 => x"81", -- $0a3b8
          41913 => x"81", -- $0a3b9
          41914 => x"81", -- $0a3ba
          41915 => x"81", -- $0a3bb
          41916 => x"80", -- $0a3bc
          41917 => x"80", -- $0a3bd
          41918 => x"80", -- $0a3be
          41919 => x"80", -- $0a3bf
          41920 => x"80", -- $0a3c0
          41921 => x"80", -- $0a3c1
          41922 => x"80", -- $0a3c2
          41923 => x"80", -- $0a3c3
          41924 => x"80", -- $0a3c4
          41925 => x"80", -- $0a3c5
          41926 => x"80", -- $0a3c6
          41927 => x"80", -- $0a3c7
          41928 => x"80", -- $0a3c8
          41929 => x"80", -- $0a3c9
          41930 => x"80", -- $0a3ca
          41931 => x"80", -- $0a3cb
          41932 => x"80", -- $0a3cc
          41933 => x"80", -- $0a3cd
          41934 => x"80", -- $0a3ce
          41935 => x"80", -- $0a3cf
          41936 => x"80", -- $0a3d0
          41937 => x"80", -- $0a3d1
          41938 => x"80", -- $0a3d2
          41939 => x"80", -- $0a3d3
          41940 => x"80", -- $0a3d4
          41941 => x"80", -- $0a3d5
          41942 => x"80", -- $0a3d6
          41943 => x"80", -- $0a3d7
          41944 => x"80", -- $0a3d8
          41945 => x"80", -- $0a3d9
          41946 => x"80", -- $0a3da
          41947 => x"80", -- $0a3db
          41948 => x"80", -- $0a3dc
          41949 => x"80", -- $0a3dd
          41950 => x"80", -- $0a3de
          41951 => x"80", -- $0a3df
          41952 => x"80", -- $0a3e0
          41953 => x"80", -- $0a3e1
          41954 => x"80", -- $0a3e2
          41955 => x"80", -- $0a3e3
          41956 => x"80", -- $0a3e4
          41957 => x"80", -- $0a3e5
          41958 => x"80", -- $0a3e6
          41959 => x"80", -- $0a3e7
          41960 => x"80", -- $0a3e8
          41961 => x"81", -- $0a3e9
          41962 => x"81", -- $0a3ea
          41963 => x"81", -- $0a3eb
          41964 => x"81", -- $0a3ec
          41965 => x"81", -- $0a3ed
          41966 => x"81", -- $0a3ee
          41967 => x"81", -- $0a3ef
          41968 => x"81", -- $0a3f0
          41969 => x"81", -- $0a3f1
          41970 => x"81", -- $0a3f2
          41971 => x"81", -- $0a3f3
          41972 => x"80", -- $0a3f4
          41973 => x"80", -- $0a3f5
          41974 => x"80", -- $0a3f6
          41975 => x"80", -- $0a3f7
          41976 => x"80", -- $0a3f8
          41977 => x"81", -- $0a3f9
          41978 => x"81", -- $0a3fa
          41979 => x"81", -- $0a3fb
          41980 => x"81", -- $0a3fc
          41981 => x"81", -- $0a3fd
          41982 => x"81", -- $0a3fe
          41983 => x"81", -- $0a3ff
          41984 => x"81", -- $0a400
          41985 => x"81", -- $0a401
          41986 => x"81", -- $0a402
          41987 => x"81", -- $0a403
          41988 => x"81", -- $0a404
          41989 => x"81", -- $0a405
          41990 => x"81", -- $0a406
          41991 => x"81", -- $0a407
          41992 => x"81", -- $0a408
          41993 => x"81", -- $0a409
          41994 => x"81", -- $0a40a
          41995 => x"81", -- $0a40b
          41996 => x"81", -- $0a40c
          41997 => x"81", -- $0a40d
          41998 => x"81", -- $0a40e
          41999 => x"80", -- $0a40f
          42000 => x"80", -- $0a410
          42001 => x"80", -- $0a411
          42002 => x"80", -- $0a412
          42003 => x"80", -- $0a413
          42004 => x"80", -- $0a414
          42005 => x"80", -- $0a415
          42006 => x"80", -- $0a416
          42007 => x"80", -- $0a417
          42008 => x"80", -- $0a418
          42009 => x"80", -- $0a419
          42010 => x"81", -- $0a41a
          42011 => x"81", -- $0a41b
          42012 => x"81", -- $0a41c
          42013 => x"81", -- $0a41d
          42014 => x"81", -- $0a41e
          42015 => x"81", -- $0a41f
          42016 => x"81", -- $0a420
          42017 => x"81", -- $0a421
          42018 => x"81", -- $0a422
          42019 => x"81", -- $0a423
          42020 => x"81", -- $0a424
          42021 => x"81", -- $0a425
          42022 => x"81", -- $0a426
          42023 => x"81", -- $0a427
          42024 => x"81", -- $0a428
          42025 => x"80", -- $0a429
          42026 => x"80", -- $0a42a
          42027 => x"80", -- $0a42b
          42028 => x"80", -- $0a42c
          42029 => x"80", -- $0a42d
          42030 => x"80", -- $0a42e
          42031 => x"80", -- $0a42f
          42032 => x"80", -- $0a430
          42033 => x"80", -- $0a431
          42034 => x"80", -- $0a432
          42035 => x"80", -- $0a433
          42036 => x"80", -- $0a434
          42037 => x"80", -- $0a435
          42038 => x"80", -- $0a436
          42039 => x"80", -- $0a437
          42040 => x"80", -- $0a438
          42041 => x"80", -- $0a439
          42042 => x"80", -- $0a43a
          42043 => x"80", -- $0a43b
          42044 => x"80", -- $0a43c
          42045 => x"80", -- $0a43d
          42046 => x"80", -- $0a43e
          42047 => x"80", -- $0a43f
          42048 => x"80", -- $0a440
          42049 => x"80", -- $0a441
          42050 => x"80", -- $0a442
          42051 => x"80", -- $0a443
          42052 => x"80", -- $0a444
          42053 => x"80", -- $0a445
          42054 => x"80", -- $0a446
          42055 => x"80", -- $0a447
          42056 => x"80", -- $0a448
          42057 => x"80", -- $0a449
          42058 => x"80", -- $0a44a
          42059 => x"80", -- $0a44b
          42060 => x"80", -- $0a44c
          42061 => x"80", -- $0a44d
          42062 => x"80", -- $0a44e
          42063 => x"80", -- $0a44f
          42064 => x"80", -- $0a450
          42065 => x"80", -- $0a451
          42066 => x"80", -- $0a452
          42067 => x"80", -- $0a453
          42068 => x"80", -- $0a454
          42069 => x"80", -- $0a455
          42070 => x"80", -- $0a456
          42071 => x"80", -- $0a457
          42072 => x"80", -- $0a458
          42073 => x"80", -- $0a459
          42074 => x"80", -- $0a45a
          42075 => x"80", -- $0a45b
          42076 => x"80", -- $0a45c
          42077 => x"80", -- $0a45d
          42078 => x"80", -- $0a45e
          42079 => x"80", -- $0a45f
          42080 => x"80", -- $0a460
          42081 => x"80", -- $0a461
          42082 => x"7f", -- $0a462
          42083 => x"7f", -- $0a463
          42084 => x"7f", -- $0a464
          42085 => x"7f", -- $0a465
          42086 => x"7f", -- $0a466
          42087 => x"7f", -- $0a467
          42088 => x"7f", -- $0a468
          42089 => x"7f", -- $0a469
          42090 => x"7f", -- $0a46a
          42091 => x"7f", -- $0a46b
          42092 => x"7f", -- $0a46c
          42093 => x"7f", -- $0a46d
          42094 => x"80", -- $0a46e
          42095 => x"80", -- $0a46f
          42096 => x"80", -- $0a470
          42097 => x"80", -- $0a471
          42098 => x"80", -- $0a472
          42099 => x"80", -- $0a473
          42100 => x"80", -- $0a474
          42101 => x"80", -- $0a475
          42102 => x"80", -- $0a476
          42103 => x"7f", -- $0a477
          42104 => x"7f", -- $0a478
          42105 => x"7f", -- $0a479
          42106 => x"7f", -- $0a47a
          42107 => x"7f", -- $0a47b
          42108 => x"7f", -- $0a47c
          42109 => x"7f", -- $0a47d
          42110 => x"7f", -- $0a47e
          42111 => x"7f", -- $0a47f
          42112 => x"7f", -- $0a480
          42113 => x"7f", -- $0a481
          42114 => x"7f", -- $0a482
          42115 => x"7f", -- $0a483
          42116 => x"7f", -- $0a484
          42117 => x"7f", -- $0a485
          42118 => x"7f", -- $0a486
          42119 => x"7f", -- $0a487
          42120 => x"7f", -- $0a488
          42121 => x"7f", -- $0a489
          42122 => x"7f", -- $0a48a
          42123 => x"7f", -- $0a48b
          42124 => x"7f", -- $0a48c
          42125 => x"7f", -- $0a48d
          42126 => x"7f", -- $0a48e
          42127 => x"7f", -- $0a48f
          42128 => x"7f", -- $0a490
          42129 => x"7f", -- $0a491
          42130 => x"7f", -- $0a492
          42131 => x"7f", -- $0a493
          42132 => x"7f", -- $0a494
          42133 => x"7f", -- $0a495
          42134 => x"7f", -- $0a496
          42135 => x"7f", -- $0a497
          42136 => x"7f", -- $0a498
          42137 => x"7f", -- $0a499
          42138 => x"7f", -- $0a49a
          42139 => x"7f", -- $0a49b
          42140 => x"7f", -- $0a49c
          42141 => x"7f", -- $0a49d
          42142 => x"7f", -- $0a49e
          42143 => x"7f", -- $0a49f
          42144 => x"7f", -- $0a4a0
          42145 => x"7f", -- $0a4a1
          42146 => x"7f", -- $0a4a2
          42147 => x"7f", -- $0a4a3
          42148 => x"80", -- $0a4a4
          42149 => x"80", -- $0a4a5
          42150 => x"80", -- $0a4a6
          42151 => x"80", -- $0a4a7
          42152 => x"80", -- $0a4a8
          42153 => x"7f", -- $0a4a9
          42154 => x"7f", -- $0a4aa
          42155 => x"7f", -- $0a4ab
          42156 => x"7f", -- $0a4ac
          42157 => x"7f", -- $0a4ad
          42158 => x"7f", -- $0a4ae
          42159 => x"7f", -- $0a4af
          42160 => x"7f", -- $0a4b0
          42161 => x"7f", -- $0a4b1
          42162 => x"7f", -- $0a4b2
          42163 => x"7f", -- $0a4b3
          42164 => x"7f", -- $0a4b4
          42165 => x"7f", -- $0a4b5
          42166 => x"7f", -- $0a4b6
          42167 => x"7f", -- $0a4b7
          42168 => x"7f", -- $0a4b8
          42169 => x"7f", -- $0a4b9
          42170 => x"7f", -- $0a4ba
          42171 => x"7f", -- $0a4bb
          42172 => x"7f", -- $0a4bc
          42173 => x"7f", -- $0a4bd
          42174 => x"7f", -- $0a4be
          42175 => x"7f", -- $0a4bf
          42176 => x"7f", -- $0a4c0
          42177 => x"7f", -- $0a4c1
          42178 => x"80", -- $0a4c2
          42179 => x"7f", -- $0a4c3
          42180 => x"7f", -- $0a4c4
          42181 => x"7f", -- $0a4c5
          42182 => x"7f", -- $0a4c6
          42183 => x"7f", -- $0a4c7
          42184 => x"7f", -- $0a4c8
          42185 => x"7f", -- $0a4c9
          42186 => x"7f", -- $0a4ca
          42187 => x"7f", -- $0a4cb
          42188 => x"7e", -- $0a4cc
          42189 => x"7e", -- $0a4cd
          42190 => x"7e", -- $0a4ce
          42191 => x"7e", -- $0a4cf
          42192 => x"7e", -- $0a4d0
          42193 => x"7e", -- $0a4d1
          42194 => x"7e", -- $0a4d2
          42195 => x"7e", -- $0a4d3
          42196 => x"7e", -- $0a4d4
          42197 => x"7f", -- $0a4d5
          42198 => x"7f", -- $0a4d6
          42199 => x"7f", -- $0a4d7
          42200 => x"7f", -- $0a4d8
          42201 => x"7f", -- $0a4d9
          42202 => x"7f", -- $0a4da
          42203 => x"7f", -- $0a4db
          42204 => x"7f", -- $0a4dc
          42205 => x"7f", -- $0a4dd
          42206 => x"7f", -- $0a4de
          42207 => x"7f", -- $0a4df
          42208 => x"7f", -- $0a4e0
          42209 => x"7f", -- $0a4e1
          42210 => x"7f", -- $0a4e2
          42211 => x"7f", -- $0a4e3
          42212 => x"7e", -- $0a4e4
          42213 => x"7e", -- $0a4e5
          42214 => x"7e", -- $0a4e6
          42215 => x"7e", -- $0a4e7
          42216 => x"7e", -- $0a4e8
          42217 => x"7e", -- $0a4e9
          42218 => x"7e", -- $0a4ea
          42219 => x"7e", -- $0a4eb
          42220 => x"7e", -- $0a4ec
          42221 => x"7e", -- $0a4ed
          42222 => x"7e", -- $0a4ee
          42223 => x"7e", -- $0a4ef
          42224 => x"7f", -- $0a4f0
          42225 => x"7f", -- $0a4f1
          42226 => x"7f", -- $0a4f2
          42227 => x"7f", -- $0a4f3
          42228 => x"7f", -- $0a4f4
          42229 => x"7f", -- $0a4f5
          42230 => x"7f", -- $0a4f6
          42231 => x"7f", -- $0a4f7
          42232 => x"7f", -- $0a4f8
          42233 => x"7f", -- $0a4f9
          42234 => x"7f", -- $0a4fa
          42235 => x"7f", -- $0a4fb
          42236 => x"7f", -- $0a4fc
          42237 => x"7f", -- $0a4fd
          42238 => x"7e", -- $0a4fe
          42239 => x"7e", -- $0a4ff
          42240 => x"7e", -- $0a500
          42241 => x"7e", -- $0a501
          42242 => x"7e", -- $0a502
          42243 => x"7e", -- $0a503
          42244 => x"7e", -- $0a504
          42245 => x"7e", -- $0a505
          42246 => x"7e", -- $0a506
          42247 => x"7e", -- $0a507
          42248 => x"7e", -- $0a508
          42249 => x"7f", -- $0a509
          42250 => x"7f", -- $0a50a
          42251 => x"7f", -- $0a50b
          42252 => x"7f", -- $0a50c
          42253 => x"7f", -- $0a50d
          42254 => x"7f", -- $0a50e
          42255 => x"7f", -- $0a50f
          42256 => x"7f", -- $0a510
          42257 => x"7f", -- $0a511
          42258 => x"7f", -- $0a512
          42259 => x"7f", -- $0a513
          42260 => x"7f", -- $0a514
          42261 => x"7f", -- $0a515
          42262 => x"7f", -- $0a516
          42263 => x"7f", -- $0a517
          42264 => x"7f", -- $0a518
          42265 => x"7f", -- $0a519
          42266 => x"7e", -- $0a51a
          42267 => x"7e", -- $0a51b
          42268 => x"7e", -- $0a51c
          42269 => x"7e", -- $0a51d
          42270 => x"7e", -- $0a51e
          42271 => x"7e", -- $0a51f
          42272 => x"7f", -- $0a520
          42273 => x"7f", -- $0a521
          42274 => x"7f", -- $0a522
          42275 => x"7f", -- $0a523
          42276 => x"7f", -- $0a524
          42277 => x"7f", -- $0a525
          42278 => x"80", -- $0a526
          42279 => x"80", -- $0a527
          42280 => x"80", -- $0a528
          42281 => x"80", -- $0a529
          42282 => x"80", -- $0a52a
          42283 => x"80", -- $0a52b
          42284 => x"80", -- $0a52c
          42285 => x"80", -- $0a52d
          42286 => x"80", -- $0a52e
          42287 => x"80", -- $0a52f
          42288 => x"80", -- $0a530
          42289 => x"7f", -- $0a531
          42290 => x"7f", -- $0a532
          42291 => x"7f", -- $0a533
          42292 => x"7f", -- $0a534
          42293 => x"7f", -- $0a535
          42294 => x"7f", -- $0a536
          42295 => x"7f", -- $0a537
          42296 => x"7f", -- $0a538
          42297 => x"7f", -- $0a539
          42298 => x"7f", -- $0a53a
          42299 => x"7f", -- $0a53b
          42300 => x"7f", -- $0a53c
          42301 => x"80", -- $0a53d
          42302 => x"80", -- $0a53e
          42303 => x"80", -- $0a53f
          42304 => x"80", -- $0a540
          42305 => x"80", -- $0a541
          42306 => x"80", -- $0a542
          42307 => x"80", -- $0a543
          42308 => x"80", -- $0a544
          42309 => x"80", -- $0a545
          42310 => x"80", -- $0a546
          42311 => x"80", -- $0a547
          42312 => x"80", -- $0a548
          42313 => x"80", -- $0a549
          42314 => x"80", -- $0a54a
          42315 => x"80", -- $0a54b
          42316 => x"7f", -- $0a54c
          42317 => x"7f", -- $0a54d
          42318 => x"7f", -- $0a54e
          42319 => x"7f", -- $0a54f
          42320 => x"7f", -- $0a550
          42321 => x"7f", -- $0a551
          42322 => x"7f", -- $0a552
          42323 => x"7f", -- $0a553
          42324 => x"7f", -- $0a554
          42325 => x"7f", -- $0a555
          42326 => x"7f", -- $0a556
          42327 => x"80", -- $0a557
          42328 => x"80", -- $0a558
          42329 => x"80", -- $0a559
          42330 => x"80", -- $0a55a
          42331 => x"80", -- $0a55b
          42332 => x"80", -- $0a55c
          42333 => x"80", -- $0a55d
          42334 => x"80", -- $0a55e
          42335 => x"80", -- $0a55f
          42336 => x"80", -- $0a560
          42337 => x"80", -- $0a561
          42338 => x"80", -- $0a562
          42339 => x"80", -- $0a563
          42340 => x"80", -- $0a564
          42341 => x"80", -- $0a565
          42342 => x"7f", -- $0a566
          42343 => x"7f", -- $0a567
          42344 => x"7f", -- $0a568
          42345 => x"7f", -- $0a569
          42346 => x"7f", -- $0a56a
          42347 => x"7f", -- $0a56b
          42348 => x"7f", -- $0a56c
          42349 => x"7f", -- $0a56d
          42350 => x"7f", -- $0a56e
          42351 => x"7f", -- $0a56f
          42352 => x"80", -- $0a570
          42353 => x"80", -- $0a571
          42354 => x"80", -- $0a572
          42355 => x"80", -- $0a573
          42356 => x"80", -- $0a574
          42357 => x"80", -- $0a575
          42358 => x"80", -- $0a576
          42359 => x"80", -- $0a577
          42360 => x"80", -- $0a578
          42361 => x"80", -- $0a579
          42362 => x"80", -- $0a57a
          42363 => x"80", -- $0a57b
          42364 => x"80", -- $0a57c
          42365 => x"80", -- $0a57d
          42366 => x"80", -- $0a57e
          42367 => x"80", -- $0a57f
          42368 => x"80", -- $0a580
          42369 => x"80", -- $0a581
          42370 => x"80", -- $0a582
          42371 => x"7f", -- $0a583
          42372 => x"7f", -- $0a584
          42373 => x"80", -- $0a585
          42374 => x"80", -- $0a586
          42375 => x"80", -- $0a587
          42376 => x"80", -- $0a588
          42377 => x"80", -- $0a589
          42378 => x"80", -- $0a58a
          42379 => x"80", -- $0a58b
          42380 => x"80", -- $0a58c
          42381 => x"80", -- $0a58d
          42382 => x"80", -- $0a58e
          42383 => x"80", -- $0a58f
          42384 => x"80", -- $0a590
          42385 => x"80", -- $0a591
          42386 => x"80", -- $0a592
          42387 => x"80", -- $0a593
          42388 => x"80", -- $0a594
          42389 => x"80", -- $0a595
          42390 => x"80", -- $0a596
          42391 => x"80", -- $0a597
          42392 => x"80", -- $0a598
          42393 => x"80", -- $0a599
          42394 => x"80", -- $0a59a
          42395 => x"80", -- $0a59b
          42396 => x"80", -- $0a59c
          42397 => x"80", -- $0a59d
          42398 => x"80", -- $0a59e
          42399 => x"80", -- $0a59f
          42400 => x"80", -- $0a5a0
          42401 => x"80", -- $0a5a1
          42402 => x"80", -- $0a5a2
          42403 => x"80", -- $0a5a3
          42404 => x"80", -- $0a5a4
          42405 => x"80", -- $0a5a5
          42406 => x"80", -- $0a5a6
          42407 => x"80", -- $0a5a7
          42408 => x"80", -- $0a5a8
          42409 => x"80", -- $0a5a9
          42410 => x"80", -- $0a5aa
          42411 => x"80", -- $0a5ab
          42412 => x"80", -- $0a5ac
          42413 => x"80", -- $0a5ad
          42414 => x"80", -- $0a5ae
          42415 => x"80", -- $0a5af
          42416 => x"80", -- $0a5b0
          42417 => x"80", -- $0a5b1
          42418 => x"80", -- $0a5b2
          42419 => x"80", -- $0a5b3
          42420 => x"80", -- $0a5b4
          42421 => x"80", -- $0a5b5
          42422 => x"80", -- $0a5b6
          42423 => x"80", -- $0a5b7
          42424 => x"80", -- $0a5b8
          42425 => x"80", -- $0a5b9
          42426 => x"80", -- $0a5ba
          42427 => x"80", -- $0a5bb
          42428 => x"80", -- $0a5bc
          42429 => x"80", -- $0a5bd
          42430 => x"80", -- $0a5be
          42431 => x"80", -- $0a5bf
          42432 => x"80", -- $0a5c0
          42433 => x"80", -- $0a5c1
          42434 => x"81", -- $0a5c2
          42435 => x"81", -- $0a5c3
          42436 => x"81", -- $0a5c4
          42437 => x"81", -- $0a5c5
          42438 => x"81", -- $0a5c6
          42439 => x"81", -- $0a5c7
          42440 => x"81", -- $0a5c8
          42441 => x"80", -- $0a5c9
          42442 => x"80", -- $0a5ca
          42443 => x"80", -- $0a5cb
          42444 => x"80", -- $0a5cc
          42445 => x"80", -- $0a5cd
          42446 => x"80", -- $0a5ce
          42447 => x"80", -- $0a5cf
          42448 => x"80", -- $0a5d0
          42449 => x"80", -- $0a5d1
          42450 => x"80", -- $0a5d2
          42451 => x"80", -- $0a5d3
          42452 => x"80", -- $0a5d4
          42453 => x"80", -- $0a5d5
          42454 => x"80", -- $0a5d6
          42455 => x"80", -- $0a5d7
          42456 => x"81", -- $0a5d8
          42457 => x"81", -- $0a5d9
          42458 => x"81", -- $0a5da
          42459 => x"81", -- $0a5db
          42460 => x"81", -- $0a5dc
          42461 => x"81", -- $0a5dd
          42462 => x"81", -- $0a5de
          42463 => x"81", -- $0a5df
          42464 => x"81", -- $0a5e0
          42465 => x"81", -- $0a5e1
          42466 => x"81", -- $0a5e2
          42467 => x"81", -- $0a5e3
          42468 => x"81", -- $0a5e4
          42469 => x"81", -- $0a5e5
          42470 => x"81", -- $0a5e6
          42471 => x"81", -- $0a5e7
          42472 => x"81", -- $0a5e8
          42473 => x"81", -- $0a5e9
          42474 => x"81", -- $0a5ea
          42475 => x"81", -- $0a5eb
          42476 => x"81", -- $0a5ec
          42477 => x"81", -- $0a5ed
          42478 => x"81", -- $0a5ee
          42479 => x"81", -- $0a5ef
          42480 => x"81", -- $0a5f0
          42481 => x"81", -- $0a5f1
          42482 => x"81", -- $0a5f2
          42483 => x"81", -- $0a5f3
          42484 => x"81", -- $0a5f4
          42485 => x"81", -- $0a5f5
          42486 => x"81", -- $0a5f6
          42487 => x"81", -- $0a5f7
          42488 => x"81", -- $0a5f8
          42489 => x"81", -- $0a5f9
          42490 => x"81", -- $0a5fa
          42491 => x"81", -- $0a5fb
          42492 => x"81", -- $0a5fc
          42493 => x"81", -- $0a5fd
          42494 => x"81", -- $0a5fe
          42495 => x"81", -- $0a5ff
          42496 => x"81", -- $0a600
          42497 => x"81", -- $0a601
          42498 => x"81", -- $0a602
          42499 => x"81", -- $0a603
          42500 => x"81", -- $0a604
          42501 => x"81", -- $0a605
          42502 => x"81", -- $0a606
          42503 => x"81", -- $0a607
          42504 => x"81", -- $0a608
          42505 => x"81", -- $0a609
          42506 => x"81", -- $0a60a
          42507 => x"81", -- $0a60b
          42508 => x"81", -- $0a60c
          42509 => x"81", -- $0a60d
          42510 => x"81", -- $0a60e
          42511 => x"81", -- $0a60f
          42512 => x"81", -- $0a610
          42513 => x"81", -- $0a611
          42514 => x"81", -- $0a612
          42515 => x"81", -- $0a613
          42516 => x"81", -- $0a614
          42517 => x"81", -- $0a615
          42518 => x"81", -- $0a616
          42519 => x"81", -- $0a617
          42520 => x"81", -- $0a618
          42521 => x"81", -- $0a619
          42522 => x"81", -- $0a61a
          42523 => x"81", -- $0a61b
          42524 => x"81", -- $0a61c
          42525 => x"81", -- $0a61d
          42526 => x"81", -- $0a61e
          42527 => x"81", -- $0a61f
          42528 => x"81", -- $0a620
          42529 => x"81", -- $0a621
          42530 => x"81", -- $0a622
          42531 => x"81", -- $0a623
          42532 => x"81", -- $0a624
          42533 => x"81", -- $0a625
          42534 => x"81", -- $0a626
          42535 => x"81", -- $0a627
          42536 => x"81", -- $0a628
          42537 => x"81", -- $0a629
          42538 => x"81", -- $0a62a
          42539 => x"81", -- $0a62b
          42540 => x"81", -- $0a62c
          42541 => x"81", -- $0a62d
          42542 => x"81", -- $0a62e
          42543 => x"81", -- $0a62f
          42544 => x"81", -- $0a630
          42545 => x"81", -- $0a631
          42546 => x"81", -- $0a632
          42547 => x"81", -- $0a633
          42548 => x"81", -- $0a634
          42549 => x"81", -- $0a635
          42550 => x"81", -- $0a636
          42551 => x"81", -- $0a637
          42552 => x"81", -- $0a638
          42553 => x"81", -- $0a639
          42554 => x"81", -- $0a63a
          42555 => x"81", -- $0a63b
          42556 => x"81", -- $0a63c
          42557 => x"81", -- $0a63d
          42558 => x"81", -- $0a63e
          42559 => x"81", -- $0a63f
          42560 => x"81", -- $0a640
          42561 => x"81", -- $0a641
          42562 => x"81", -- $0a642
          42563 => x"81", -- $0a643
          42564 => x"81", -- $0a644
          42565 => x"81", -- $0a645
          42566 => x"81", -- $0a646
          42567 => x"81", -- $0a647
          42568 => x"81", -- $0a648
          42569 => x"81", -- $0a649
          42570 => x"81", -- $0a64a
          42571 => x"81", -- $0a64b
          42572 => x"81", -- $0a64c
          42573 => x"81", -- $0a64d
          42574 => x"81", -- $0a64e
          42575 => x"81", -- $0a64f
          42576 => x"81", -- $0a650
          42577 => x"81", -- $0a651
          42578 => x"81", -- $0a652
          42579 => x"81", -- $0a653
          42580 => x"81", -- $0a654
          42581 => x"81", -- $0a655
          42582 => x"81", -- $0a656
          42583 => x"81", -- $0a657
          42584 => x"81", -- $0a658
          42585 => x"81", -- $0a659
          42586 => x"81", -- $0a65a
          42587 => x"81", -- $0a65b
          42588 => x"81", -- $0a65c
          42589 => x"81", -- $0a65d
          42590 => x"81", -- $0a65e
          42591 => x"81", -- $0a65f
          42592 => x"81", -- $0a660
          42593 => x"81", -- $0a661
          42594 => x"81", -- $0a662
          42595 => x"81", -- $0a663
          42596 => x"81", -- $0a664
          42597 => x"81", -- $0a665
          42598 => x"81", -- $0a666
          42599 => x"81", -- $0a667
          42600 => x"81", -- $0a668
          42601 => x"81", -- $0a669
          42602 => x"81", -- $0a66a
          42603 => x"81", -- $0a66b
          42604 => x"81", -- $0a66c
          42605 => x"81", -- $0a66d
          42606 => x"81", -- $0a66e
          42607 => x"81", -- $0a66f
          42608 => x"81", -- $0a670
          42609 => x"81", -- $0a671
          42610 => x"81", -- $0a672
          42611 => x"81", -- $0a673
          42612 => x"81", -- $0a674
          42613 => x"81", -- $0a675
          42614 => x"81", -- $0a676
          42615 => x"81", -- $0a677
          42616 => x"81", -- $0a678
          42617 => x"81", -- $0a679
          42618 => x"81", -- $0a67a
          42619 => x"81", -- $0a67b
          42620 => x"81", -- $0a67c
          42621 => x"81", -- $0a67d
          42622 => x"81", -- $0a67e
          42623 => x"81", -- $0a67f
          42624 => x"81", -- $0a680
          42625 => x"81", -- $0a681
          42626 => x"81", -- $0a682
          42627 => x"81", -- $0a683
          42628 => x"81", -- $0a684
          42629 => x"81", -- $0a685
          42630 => x"81", -- $0a686
          42631 => x"81", -- $0a687
          42632 => x"81", -- $0a688
          42633 => x"81", -- $0a689
          42634 => x"81", -- $0a68a
          42635 => x"81", -- $0a68b
          42636 => x"81", -- $0a68c
          42637 => x"81", -- $0a68d
          42638 => x"81", -- $0a68e
          42639 => x"81", -- $0a68f
          42640 => x"81", -- $0a690
          42641 => x"81", -- $0a691
          42642 => x"81", -- $0a692
          42643 => x"81", -- $0a693
          42644 => x"81", -- $0a694
          42645 => x"81", -- $0a695
          42646 => x"81", -- $0a696
          42647 => x"81", -- $0a697
          42648 => x"81", -- $0a698
          42649 => x"81", -- $0a699
          42650 => x"81", -- $0a69a
          42651 => x"81", -- $0a69b
          42652 => x"81", -- $0a69c
          42653 => x"81", -- $0a69d
          42654 => x"81", -- $0a69e
          42655 => x"81", -- $0a69f
          42656 => x"81", -- $0a6a0
          42657 => x"81", -- $0a6a1
          42658 => x"81", -- $0a6a2
          42659 => x"81", -- $0a6a3
          42660 => x"81", -- $0a6a4
          42661 => x"81", -- $0a6a5
          42662 => x"81", -- $0a6a6
          42663 => x"81", -- $0a6a7
          42664 => x"81", -- $0a6a8
          42665 => x"81", -- $0a6a9
          42666 => x"81", -- $0a6aa
          42667 => x"81", -- $0a6ab
          42668 => x"81", -- $0a6ac
          42669 => x"81", -- $0a6ad
          42670 => x"81", -- $0a6ae
          42671 => x"81", -- $0a6af
          42672 => x"81", -- $0a6b0
          42673 => x"81", -- $0a6b1
          42674 => x"81", -- $0a6b2
          42675 => x"81", -- $0a6b3
          42676 => x"81", -- $0a6b4
          42677 => x"81", -- $0a6b5
          42678 => x"81", -- $0a6b6
          42679 => x"81", -- $0a6b7
          42680 => x"81", -- $0a6b8
          42681 => x"81", -- $0a6b9
          42682 => x"81", -- $0a6ba
          42683 => x"81", -- $0a6bb
          42684 => x"81", -- $0a6bc
          42685 => x"81", -- $0a6bd
          42686 => x"81", -- $0a6be
          42687 => x"80", -- $0a6bf
          42688 => x"80", -- $0a6c0
          42689 => x"80", -- $0a6c1
          42690 => x"80", -- $0a6c2
          42691 => x"80", -- $0a6c3
          42692 => x"80", -- $0a6c4
          42693 => x"80", -- $0a6c5
          42694 => x"80", -- $0a6c6
          42695 => x"80", -- $0a6c7
          42696 => x"80", -- $0a6c8
          42697 => x"80", -- $0a6c9
          42698 => x"80", -- $0a6ca
          42699 => x"80", -- $0a6cb
          42700 => x"80", -- $0a6cc
          42701 => x"80", -- $0a6cd
          42702 => x"80", -- $0a6ce
          42703 => x"80", -- $0a6cf
          42704 => x"80", -- $0a6d0
          42705 => x"80", -- $0a6d1
          42706 => x"80", -- $0a6d2
          42707 => x"81", -- $0a6d3
          42708 => x"80", -- $0a6d4
          42709 => x"81", -- $0a6d5
          42710 => x"80", -- $0a6d6
          42711 => x"80", -- $0a6d7
          42712 => x"80", -- $0a6d8
          42713 => x"80", -- $0a6d9
          42714 => x"80", -- $0a6da
          42715 => x"80", -- $0a6db
          42716 => x"80", -- $0a6dc
          42717 => x"80", -- $0a6dd
          42718 => x"80", -- $0a6de
          42719 => x"80", -- $0a6df
          42720 => x"80", -- $0a6e0
          42721 => x"80", -- $0a6e1
          42722 => x"80", -- $0a6e2
          42723 => x"80", -- $0a6e3
          42724 => x"80", -- $0a6e4
          42725 => x"80", -- $0a6e5
          42726 => x"80", -- $0a6e6
          42727 => x"80", -- $0a6e7
          42728 => x"80", -- $0a6e8
          42729 => x"80", -- $0a6e9
          42730 => x"80", -- $0a6ea
          42731 => x"80", -- $0a6eb
          42732 => x"80", -- $0a6ec
          42733 => x"80", -- $0a6ed
          42734 => x"80", -- $0a6ee
          42735 => x"80", -- $0a6ef
          42736 => x"80", -- $0a6f0
          42737 => x"80", -- $0a6f1
          42738 => x"80", -- $0a6f2
          42739 => x"80", -- $0a6f3
          42740 => x"80", -- $0a6f4
          42741 => x"80", -- $0a6f5
          42742 => x"80", -- $0a6f6
          42743 => x"80", -- $0a6f7
          42744 => x"80", -- $0a6f8
          42745 => x"80", -- $0a6f9
          42746 => x"80", -- $0a6fa
          42747 => x"80", -- $0a6fb
          42748 => x"80", -- $0a6fc
          42749 => x"80", -- $0a6fd
          42750 => x"80", -- $0a6fe
          42751 => x"80", -- $0a6ff
          42752 => x"80", -- $0a700
          42753 => x"80", -- $0a701
          42754 => x"80", -- $0a702
          42755 => x"80", -- $0a703
          42756 => x"80", -- $0a704
          42757 => x"80", -- $0a705
          42758 => x"80", -- $0a706
          42759 => x"80", -- $0a707
          42760 => x"80", -- $0a708
          42761 => x"80", -- $0a709
          42762 => x"80", -- $0a70a
          42763 => x"80", -- $0a70b
          42764 => x"80", -- $0a70c
          42765 => x"80", -- $0a70d
          42766 => x"80", -- $0a70e
          42767 => x"80", -- $0a70f
          42768 => x"80", -- $0a710
          42769 => x"80", -- $0a711
          42770 => x"7f", -- $0a712
          42771 => x"7f", -- $0a713
          42772 => x"7f", -- $0a714
          42773 => x"80", -- $0a715
          42774 => x"7f", -- $0a716
          42775 => x"7f", -- $0a717
          42776 => x"80", -- $0a718
          42777 => x"80", -- $0a719
          42778 => x"80", -- $0a71a
          42779 => x"80", -- $0a71b
          42780 => x"80", -- $0a71c
          42781 => x"80", -- $0a71d
          42782 => x"80", -- $0a71e
          42783 => x"80", -- $0a71f
          42784 => x"80", -- $0a720
          42785 => x"80", -- $0a721
          42786 => x"80", -- $0a722
          42787 => x"80", -- $0a723
          42788 => x"80", -- $0a724
          42789 => x"80", -- $0a725
          42790 => x"80", -- $0a726
          42791 => x"80", -- $0a727
          42792 => x"80", -- $0a728
          42793 => x"80", -- $0a729
          42794 => x"7f", -- $0a72a
          42795 => x"7f", -- $0a72b
          42796 => x"7f", -- $0a72c
          42797 => x"7f", -- $0a72d
          42798 => x"7f", -- $0a72e
          42799 => x"7f", -- $0a72f
          42800 => x"7f", -- $0a730
          42801 => x"7f", -- $0a731
          42802 => x"7f", -- $0a732
          42803 => x"7f", -- $0a733
          42804 => x"80", -- $0a734
          42805 => x"80", -- $0a735
          42806 => x"7f", -- $0a736
          42807 => x"80", -- $0a737
          42808 => x"80", -- $0a738
          42809 => x"80", -- $0a739
          42810 => x"80", -- $0a73a
          42811 => x"80", -- $0a73b
          42812 => x"80", -- $0a73c
          42813 => x"80", -- $0a73d
          42814 => x"80", -- $0a73e
          42815 => x"80", -- $0a73f
          42816 => x"80", -- $0a740
          42817 => x"80", -- $0a741
          42818 => x"7f", -- $0a742
          42819 => x"7f", -- $0a743
          42820 => x"7f", -- $0a744
          42821 => x"7f", -- $0a745
          42822 => x"7f", -- $0a746
          42823 => x"7f", -- $0a747
          42824 => x"7f", -- $0a748
          42825 => x"7f", -- $0a749
          42826 => x"7f", -- $0a74a
          42827 => x"7f", -- $0a74b
          42828 => x"7f", -- $0a74c
          42829 => x"7f", -- $0a74d
          42830 => x"7f", -- $0a74e
          42831 => x"7f", -- $0a74f
          42832 => x"7f", -- $0a750
          42833 => x"7f", -- $0a751
          42834 => x"7f", -- $0a752
          42835 => x"80", -- $0a753
          42836 => x"80", -- $0a754
          42837 => x"80", -- $0a755
          42838 => x"80", -- $0a756
          42839 => x"80", -- $0a757
          42840 => x"80", -- $0a758
          42841 => x"80", -- $0a759
          42842 => x"80", -- $0a75a
          42843 => x"80", -- $0a75b
          42844 => x"7f", -- $0a75c
          42845 => x"7f", -- $0a75d
          42846 => x"7f", -- $0a75e
          42847 => x"7f", -- $0a75f
          42848 => x"7f", -- $0a760
          42849 => x"7f", -- $0a761
          42850 => x"7f", -- $0a762
          42851 => x"7f", -- $0a763
          42852 => x"7f", -- $0a764
          42853 => x"7f", -- $0a765
          42854 => x"7f", -- $0a766
          42855 => x"7f", -- $0a767
          42856 => x"7f", -- $0a768
          42857 => x"7f", -- $0a769
          42858 => x"7f", -- $0a76a
          42859 => x"7f", -- $0a76b
          42860 => x"7f", -- $0a76c
          42861 => x"7f", -- $0a76d
          42862 => x"80", -- $0a76e
          42863 => x"80", -- $0a76f
          42864 => x"80", -- $0a770
          42865 => x"80", -- $0a771
          42866 => x"80", -- $0a772
          42867 => x"80", -- $0a773
          42868 => x"80", -- $0a774
          42869 => x"80", -- $0a775
          42870 => x"80", -- $0a776
          42871 => x"80", -- $0a777
          42872 => x"7f", -- $0a778
          42873 => x"7f", -- $0a779
          42874 => x"7f", -- $0a77a
          42875 => x"7f", -- $0a77b
          42876 => x"7f", -- $0a77c
          42877 => x"7f", -- $0a77d
          42878 => x"7f", -- $0a77e
          42879 => x"7f", -- $0a77f
          42880 => x"7f", -- $0a780
          42881 => x"7f", -- $0a781
          42882 => x"7f", -- $0a782
          42883 => x"7f", -- $0a783
          42884 => x"7f", -- $0a784
          42885 => x"7f", -- $0a785
          42886 => x"7f", -- $0a786
          42887 => x"80", -- $0a787
          42888 => x"80", -- $0a788
          42889 => x"80", -- $0a789
          42890 => x"80", -- $0a78a
          42891 => x"80", -- $0a78b
          42892 => x"80", -- $0a78c
          42893 => x"80", -- $0a78d
          42894 => x"80", -- $0a78e
          42895 => x"80", -- $0a78f
          42896 => x"80", -- $0a790
          42897 => x"80", -- $0a791
          42898 => x"80", -- $0a792
          42899 => x"7f", -- $0a793
          42900 => x"7f", -- $0a794
          42901 => x"7f", -- $0a795
          42902 => x"7f", -- $0a796
          42903 => x"7f", -- $0a797
          42904 => x"7f", -- $0a798
          42905 => x"7f", -- $0a799
          42906 => x"7f", -- $0a79a
          42907 => x"7f", -- $0a79b
          42908 => x"7f", -- $0a79c
          42909 => x"7f", -- $0a79d
          42910 => x"7f", -- $0a79e
          42911 => x"7f", -- $0a79f
          42912 => x"80", -- $0a7a0
          42913 => x"80", -- $0a7a1
          42914 => x"80", -- $0a7a2
          42915 => x"80", -- $0a7a3
          42916 => x"80", -- $0a7a4
          42917 => x"80", -- $0a7a5
          42918 => x"80", -- $0a7a6
          42919 => x"80", -- $0a7a7
          42920 => x"80", -- $0a7a8
          42921 => x"80", -- $0a7a9
          42922 => x"80", -- $0a7aa
          42923 => x"80", -- $0a7ab
          42924 => x"80", -- $0a7ac
          42925 => x"7f", -- $0a7ad
          42926 => x"7f", -- $0a7ae
          42927 => x"7f", -- $0a7af
          42928 => x"7f", -- $0a7b0
          42929 => x"7f", -- $0a7b1
          42930 => x"7f", -- $0a7b2
          42931 => x"7f", -- $0a7b3
          42932 => x"7f", -- $0a7b4
          42933 => x"7f", -- $0a7b5
          42934 => x"7f", -- $0a7b6
          42935 => x"7f", -- $0a7b7
          42936 => x"7f", -- $0a7b8
          42937 => x"7f", -- $0a7b9
          42938 => x"7f", -- $0a7ba
          42939 => x"7f", -- $0a7bb
          42940 => x"7f", -- $0a7bc
          42941 => x"7f", -- $0a7bd
          42942 => x"80", -- $0a7be
          42943 => x"80", -- $0a7bf
          42944 => x"80", -- $0a7c0
          42945 => x"80", -- $0a7c1
          42946 => x"80", -- $0a7c2
          42947 => x"80", -- $0a7c3
          42948 => x"80", -- $0a7c4
          42949 => x"80", -- $0a7c5
          42950 => x"80", -- $0a7c6
          42951 => x"80", -- $0a7c7
          42952 => x"7f", -- $0a7c8
          42953 => x"7f", -- $0a7c9
          42954 => x"7f", -- $0a7ca
          42955 => x"7f", -- $0a7cb
          42956 => x"7f", -- $0a7cc
          42957 => x"7f", -- $0a7cd
          42958 => x"7f", -- $0a7ce
          42959 => x"7f", -- $0a7cf
          42960 => x"7f", -- $0a7d0
          42961 => x"7f", -- $0a7d1
          42962 => x"7f", -- $0a7d2
          42963 => x"7f", -- $0a7d3
          42964 => x"7f", -- $0a7d4
          42965 => x"7f", -- $0a7d5
          42966 => x"7f", -- $0a7d6
          42967 => x"7f", -- $0a7d7
          42968 => x"7f", -- $0a7d8
          42969 => x"7f", -- $0a7d9
          42970 => x"80", -- $0a7da
          42971 => x"7f", -- $0a7db
          42972 => x"7f", -- $0a7dc
          42973 => x"7f", -- $0a7dd
          42974 => x"7f", -- $0a7de
          42975 => x"7f", -- $0a7df
          42976 => x"7f", -- $0a7e0
          42977 => x"7f", -- $0a7e1
          42978 => x"7f", -- $0a7e2
          42979 => x"7f", -- $0a7e3
          42980 => x"7e", -- $0a7e4
          42981 => x"7e", -- $0a7e5
          42982 => x"7e", -- $0a7e6
          42983 => x"7e", -- $0a7e7
          42984 => x"7e", -- $0a7e8
          42985 => x"7e", -- $0a7e9
          42986 => x"7e", -- $0a7ea
          42987 => x"7e", -- $0a7eb
          42988 => x"7e", -- $0a7ec
          42989 => x"7e", -- $0a7ed
          42990 => x"7e", -- $0a7ee
          42991 => x"7e", -- $0a7ef
          42992 => x"7e", -- $0a7f0
          42993 => x"7f", -- $0a7f1
          42994 => x"7f", -- $0a7f2
          42995 => x"7f", -- $0a7f3
          42996 => x"7f", -- $0a7f4
          42997 => x"7f", -- $0a7f5
          42998 => x"7f", -- $0a7f6
          42999 => x"7f", -- $0a7f7
          43000 => x"7f", -- $0a7f8
          43001 => x"7f", -- $0a7f9
          43002 => x"7f", -- $0a7fa
          43003 => x"7f", -- $0a7fb
          43004 => x"7f", -- $0a7fc
          43005 => x"7e", -- $0a7fd
          43006 => x"7e", -- $0a7fe
          43007 => x"7e", -- $0a7ff
          43008 => x"7f", -- $0a800
          43009 => x"7e", -- $0a801
          43010 => x"7e", -- $0a802
          43011 => x"7e", -- $0a803
          43012 => x"7f", -- $0a804
          43013 => x"7e", -- $0a805
          43014 => x"7e", -- $0a806
          43015 => x"7e", -- $0a807
          43016 => x"7f", -- $0a808
          43017 => x"7f", -- $0a809
          43018 => x"7f", -- $0a80a
          43019 => x"7f", -- $0a80b
          43020 => x"7f", -- $0a80c
          43021 => x"7f", -- $0a80d
          43022 => x"7f", -- $0a80e
          43023 => x"7f", -- $0a80f
          43024 => x"7f", -- $0a810
          43025 => x"7f", -- $0a811
          43026 => x"7f", -- $0a812
          43027 => x"7f", -- $0a813
          43028 => x"7f", -- $0a814
          43029 => x"7f", -- $0a815
          43030 => x"7f", -- $0a816
          43031 => x"7f", -- $0a817
          43032 => x"7f", -- $0a818
          43033 => x"7f", -- $0a819
          43034 => x"7f", -- $0a81a
          43035 => x"7f", -- $0a81b
          43036 => x"7f", -- $0a81c
          43037 => x"7f", -- $0a81d
          43038 => x"7f", -- $0a81e
          43039 => x"7f", -- $0a81f
          43040 => x"7f", -- $0a820
          43041 => x"7f", -- $0a821
          43042 => x"7f", -- $0a822
          43043 => x"7f", -- $0a823
          43044 => x"80", -- $0a824
          43045 => x"80", -- $0a825
          43046 => x"80", -- $0a826
          43047 => x"80", -- $0a827
          43048 => x"80", -- $0a828
          43049 => x"80", -- $0a829
          43050 => x"80", -- $0a82a
          43051 => x"80", -- $0a82b
          43052 => x"80", -- $0a82c
          43053 => x"80", -- $0a82d
          43054 => x"80", -- $0a82e
          43055 => x"80", -- $0a82f
          43056 => x"80", -- $0a830
          43057 => x"80", -- $0a831
          43058 => x"80", -- $0a832
          43059 => x"80", -- $0a833
          43060 => x"80", -- $0a834
          43061 => x"80", -- $0a835
          43062 => x"80", -- $0a836
          43063 => x"80", -- $0a837
          43064 => x"80", -- $0a838
          43065 => x"80", -- $0a839
          43066 => x"80", -- $0a83a
          43067 => x"80", -- $0a83b
          43068 => x"80", -- $0a83c
          43069 => x"80", -- $0a83d
          43070 => x"80", -- $0a83e
          43071 => x"80", -- $0a83f
          43072 => x"80", -- $0a840
          43073 => x"80", -- $0a841
          43074 => x"80", -- $0a842
          43075 => x"80", -- $0a843
          43076 => x"80", -- $0a844
          43077 => x"80", -- $0a845
          43078 => x"80", -- $0a846
          43079 => x"80", -- $0a847
          43080 => x"80", -- $0a848
          43081 => x"80", -- $0a849
          43082 => x"80", -- $0a84a
          43083 => x"80", -- $0a84b
          43084 => x"80", -- $0a84c
          43085 => x"80", -- $0a84d
          43086 => x"80", -- $0a84e
          43087 => x"80", -- $0a84f
          43088 => x"80", -- $0a850
          43089 => x"80", -- $0a851
          43090 => x"80", -- $0a852
          43091 => x"80", -- $0a853
          43092 => x"80", -- $0a854
          43093 => x"80", -- $0a855
          43094 => x"80", -- $0a856
          43095 => x"80", -- $0a857
          43096 => x"80", -- $0a858
          43097 => x"80", -- $0a859
          43098 => x"80", -- $0a85a
          43099 => x"80", -- $0a85b
          43100 => x"80", -- $0a85c
          43101 => x"80", -- $0a85d
          43102 => x"80", -- $0a85e
          43103 => x"80", -- $0a85f
          43104 => x"80", -- $0a860
          43105 => x"80", -- $0a861
          43106 => x"80", -- $0a862
          43107 => x"80", -- $0a863
          43108 => x"80", -- $0a864
          43109 => x"80", -- $0a865
          43110 => x"80", -- $0a866
          43111 => x"80", -- $0a867
          43112 => x"80", -- $0a868
          43113 => x"80", -- $0a869
          43114 => x"80", -- $0a86a
          43115 => x"80", -- $0a86b
          43116 => x"80", -- $0a86c
          43117 => x"80", -- $0a86d
          43118 => x"80", -- $0a86e
          43119 => x"80", -- $0a86f
          43120 => x"80", -- $0a870
          43121 => x"80", -- $0a871
          43122 => x"80", -- $0a872
          43123 => x"80", -- $0a873
          43124 => x"80", -- $0a874
          43125 => x"80", -- $0a875
          43126 => x"81", -- $0a876
          43127 => x"81", -- $0a877
          43128 => x"81", -- $0a878
          43129 => x"81", -- $0a879
          43130 => x"81", -- $0a87a
          43131 => x"80", -- $0a87b
          43132 => x"80", -- $0a87c
          43133 => x"80", -- $0a87d
          43134 => x"80", -- $0a87e
          43135 => x"80", -- $0a87f
          43136 => x"80", -- $0a880
          43137 => x"80", -- $0a881
          43138 => x"80", -- $0a882
          43139 => x"80", -- $0a883
          43140 => x"80", -- $0a884
          43141 => x"80", -- $0a885
          43142 => x"80", -- $0a886
          43143 => x"80", -- $0a887
          43144 => x"80", -- $0a888
          43145 => x"80", -- $0a889
          43146 => x"80", -- $0a88a
          43147 => x"80", -- $0a88b
          43148 => x"81", -- $0a88c
          43149 => x"81", -- $0a88d
          43150 => x"81", -- $0a88e
          43151 => x"81", -- $0a88f
          43152 => x"81", -- $0a890
          43153 => x"81", -- $0a891
          43154 => x"81", -- $0a892
          43155 => x"81", -- $0a893
          43156 => x"81", -- $0a894
          43157 => x"81", -- $0a895
          43158 => x"81", -- $0a896
          43159 => x"81", -- $0a897
          43160 => x"80", -- $0a898
          43161 => x"80", -- $0a899
          43162 => x"80", -- $0a89a
          43163 => x"80", -- $0a89b
          43164 => x"80", -- $0a89c
          43165 => x"80", -- $0a89d
          43166 => x"80", -- $0a89e
          43167 => x"80", -- $0a89f
          43168 => x"80", -- $0a8a0
          43169 => x"80", -- $0a8a1
          43170 => x"80", -- $0a8a2
          43171 => x"80", -- $0a8a3
          43172 => x"80", -- $0a8a4
          43173 => x"80", -- $0a8a5
          43174 => x"80", -- $0a8a6
          43175 => x"80", -- $0a8a7
          43176 => x"80", -- $0a8a8
          43177 => x"80", -- $0a8a9
          43178 => x"80", -- $0a8aa
          43179 => x"81", -- $0a8ab
          43180 => x"81", -- $0a8ac
          43181 => x"81", -- $0a8ad
          43182 => x"81", -- $0a8ae
          43183 => x"81", -- $0a8af
          43184 => x"80", -- $0a8b0
          43185 => x"80", -- $0a8b1
          43186 => x"80", -- $0a8b2
          43187 => x"80", -- $0a8b3
          43188 => x"80", -- $0a8b4
          43189 => x"80", -- $0a8b5
          43190 => x"80", -- $0a8b6
          43191 => x"80", -- $0a8b7
          43192 => x"80", -- $0a8b8
          43193 => x"80", -- $0a8b9
          43194 => x"80", -- $0a8ba
          43195 => x"80", -- $0a8bb
          43196 => x"80", -- $0a8bc
          43197 => x"80", -- $0a8bd
          43198 => x"80", -- $0a8be
          43199 => x"80", -- $0a8bf
          43200 => x"80", -- $0a8c0
          43201 => x"80", -- $0a8c1
          43202 => x"80", -- $0a8c2
          43203 => x"81", -- $0a8c3
          43204 => x"81", -- $0a8c4
          43205 => x"81", -- $0a8c5
          43206 => x"81", -- $0a8c6
          43207 => x"81", -- $0a8c7
          43208 => x"81", -- $0a8c8
          43209 => x"81", -- $0a8c9
          43210 => x"81", -- $0a8ca
          43211 => x"81", -- $0a8cb
          43212 => x"81", -- $0a8cc
          43213 => x"80", -- $0a8cd
          43214 => x"80", -- $0a8ce
          43215 => x"80", -- $0a8cf
          43216 => x"80", -- $0a8d0
          43217 => x"80", -- $0a8d1
          43218 => x"80", -- $0a8d2
          43219 => x"80", -- $0a8d3
          43220 => x"80", -- $0a8d4
          43221 => x"80", -- $0a8d5
          43222 => x"80", -- $0a8d6
          43223 => x"80", -- $0a8d7
          43224 => x"80", -- $0a8d8
          43225 => x"80", -- $0a8d9
          43226 => x"80", -- $0a8da
          43227 => x"80", -- $0a8db
          43228 => x"80", -- $0a8dc
          43229 => x"80", -- $0a8dd
          43230 => x"80", -- $0a8de
          43231 => x"81", -- $0a8df
          43232 => x"81", -- $0a8e0
          43233 => x"81", -- $0a8e1
          43234 => x"81", -- $0a8e2
          43235 => x"81", -- $0a8e3
          43236 => x"81", -- $0a8e4
          43237 => x"81", -- $0a8e5
          43238 => x"81", -- $0a8e6
          43239 => x"81", -- $0a8e7
          43240 => x"81", -- $0a8e8
          43241 => x"81", -- $0a8e9
          43242 => x"81", -- $0a8ea
          43243 => x"81", -- $0a8eb
          43244 => x"81", -- $0a8ec
          43245 => x"81", -- $0a8ed
          43246 => x"81", -- $0a8ee
          43247 => x"80", -- $0a8ef
          43248 => x"80", -- $0a8f0
          43249 => x"80", -- $0a8f1
          43250 => x"81", -- $0a8f2
          43251 => x"81", -- $0a8f3
          43252 => x"80", -- $0a8f4
          43253 => x"81", -- $0a8f5
          43254 => x"81", -- $0a8f6
          43255 => x"81", -- $0a8f7
          43256 => x"81", -- $0a8f8
          43257 => x"81", -- $0a8f9
          43258 => x"81", -- $0a8fa
          43259 => x"81", -- $0a8fb
          43260 => x"81", -- $0a8fc
          43261 => x"81", -- $0a8fd
          43262 => x"81", -- $0a8fe
          43263 => x"81", -- $0a8ff
          43264 => x"81", -- $0a900
          43265 => x"81", -- $0a901
          43266 => x"81", -- $0a902
          43267 => x"81", -- $0a903
          43268 => x"81", -- $0a904
          43269 => x"81", -- $0a905
          43270 => x"81", -- $0a906
          43271 => x"81", -- $0a907
          43272 => x"81", -- $0a908
          43273 => x"81", -- $0a909
          43274 => x"81", -- $0a90a
          43275 => x"81", -- $0a90b
          43276 => x"81", -- $0a90c
          43277 => x"81", -- $0a90d
          43278 => x"81", -- $0a90e
          43279 => x"81", -- $0a90f
          43280 => x"81", -- $0a910
          43281 => x"81", -- $0a911
          43282 => x"81", -- $0a912
          43283 => x"81", -- $0a913
          43284 => x"81", -- $0a914
          43285 => x"81", -- $0a915
          43286 => x"81", -- $0a916
          43287 => x"81", -- $0a917
          43288 => x"81", -- $0a918
          43289 => x"81", -- $0a919
          43290 => x"81", -- $0a91a
          43291 => x"81", -- $0a91b
          43292 => x"81", -- $0a91c
          43293 => x"81", -- $0a91d
          43294 => x"81", -- $0a91e
          43295 => x"81", -- $0a91f
          43296 => x"81", -- $0a920
          43297 => x"81", -- $0a921
          43298 => x"81", -- $0a922
          43299 => x"81", -- $0a923
          43300 => x"81", -- $0a924
          43301 => x"81", -- $0a925
          43302 => x"81", -- $0a926
          43303 => x"81", -- $0a927
          43304 => x"81", -- $0a928
          43305 => x"81", -- $0a929
          43306 => x"81", -- $0a92a
          43307 => x"81", -- $0a92b
          43308 => x"81", -- $0a92c
          43309 => x"81", -- $0a92d
          43310 => x"81", -- $0a92e
          43311 => x"81", -- $0a92f
          43312 => x"81", -- $0a930
          43313 => x"81", -- $0a931
          43314 => x"81", -- $0a932
          43315 => x"81", -- $0a933
          43316 => x"81", -- $0a934
          43317 => x"81", -- $0a935
          43318 => x"81", -- $0a936
          43319 => x"81", -- $0a937
          43320 => x"81", -- $0a938
          43321 => x"81", -- $0a939
          43322 => x"81", -- $0a93a
          43323 => x"81", -- $0a93b
          43324 => x"81", -- $0a93c
          43325 => x"81", -- $0a93d
          43326 => x"81", -- $0a93e
          43327 => x"81", -- $0a93f
          43328 => x"81", -- $0a940
          43329 => x"81", -- $0a941
          43330 => x"81", -- $0a942
          43331 => x"81", -- $0a943
          43332 => x"81", -- $0a944
          43333 => x"81", -- $0a945
          43334 => x"81", -- $0a946
          43335 => x"81", -- $0a947
          43336 => x"81", -- $0a948
          43337 => x"81", -- $0a949
          43338 => x"81", -- $0a94a
          43339 => x"81", -- $0a94b
          43340 => x"81", -- $0a94c
          43341 => x"81", -- $0a94d
          43342 => x"81", -- $0a94e
          43343 => x"81", -- $0a94f
          43344 => x"81", -- $0a950
          43345 => x"81", -- $0a951
          43346 => x"81", -- $0a952
          43347 => x"81", -- $0a953
          43348 => x"81", -- $0a954
          43349 => x"81", -- $0a955
          43350 => x"81", -- $0a956
          43351 => x"81", -- $0a957
          43352 => x"81", -- $0a958
          43353 => x"80", -- $0a959
          43354 => x"81", -- $0a95a
          43355 => x"81", -- $0a95b
          43356 => x"81", -- $0a95c
          43357 => x"81", -- $0a95d
          43358 => x"81", -- $0a95e
          43359 => x"81", -- $0a95f
          43360 => x"81", -- $0a960
          43361 => x"81", -- $0a961
          43362 => x"81", -- $0a962
          43363 => x"81", -- $0a963
          43364 => x"81", -- $0a964
          43365 => x"81", -- $0a965
          43366 => x"81", -- $0a966
          43367 => x"81", -- $0a967
          43368 => x"81", -- $0a968
          43369 => x"80", -- $0a969
          43370 => x"80", -- $0a96a
          43371 => x"80", -- $0a96b
          43372 => x"80", -- $0a96c
          43373 => x"80", -- $0a96d
          43374 => x"81", -- $0a96e
          43375 => x"81", -- $0a96f
          43376 => x"80", -- $0a970
          43377 => x"80", -- $0a971
          43378 => x"80", -- $0a972
          43379 => x"80", -- $0a973
          43380 => x"80", -- $0a974
          43381 => x"80", -- $0a975
          43382 => x"80", -- $0a976
          43383 => x"80", -- $0a977
          43384 => x"80", -- $0a978
          43385 => x"80", -- $0a979
          43386 => x"80", -- $0a97a
          43387 => x"80", -- $0a97b
          43388 => x"80", -- $0a97c
          43389 => x"80", -- $0a97d
          43390 => x"80", -- $0a97e
          43391 => x"80", -- $0a97f
          43392 => x"80", -- $0a980
          43393 => x"80", -- $0a981
          43394 => x"80", -- $0a982
          43395 => x"80", -- $0a983
          43396 => x"80", -- $0a984
          43397 => x"80", -- $0a985
          43398 => x"80", -- $0a986
          43399 => x"80", -- $0a987
          43400 => x"80", -- $0a988
          43401 => x"80", -- $0a989
          43402 => x"80", -- $0a98a
          43403 => x"80", -- $0a98b
          43404 => x"80", -- $0a98c
          43405 => x"80", -- $0a98d
          43406 => x"80", -- $0a98e
          43407 => x"80", -- $0a98f
          43408 => x"80", -- $0a990
          43409 => x"80", -- $0a991
          43410 => x"80", -- $0a992
          43411 => x"80", -- $0a993
          43412 => x"80", -- $0a994
          43413 => x"80", -- $0a995
          43414 => x"80", -- $0a996
          43415 => x"80", -- $0a997
          43416 => x"80", -- $0a998
          43417 => x"80", -- $0a999
          43418 => x"80", -- $0a99a
          43419 => x"80", -- $0a99b
          43420 => x"80", -- $0a99c
          43421 => x"80", -- $0a99d
          43422 => x"80", -- $0a99e
          43423 => x"80", -- $0a99f
          43424 => x"80", -- $0a9a0
          43425 => x"80", -- $0a9a1
          43426 => x"80", -- $0a9a2
          43427 => x"80", -- $0a9a3
          43428 => x"80", -- $0a9a4
          43429 => x"80", -- $0a9a5
          43430 => x"80", -- $0a9a6
          43431 => x"80", -- $0a9a7
          43432 => x"80", -- $0a9a8
          43433 => x"80", -- $0a9a9
          43434 => x"80", -- $0a9aa
          43435 => x"80", -- $0a9ab
          43436 => x"80", -- $0a9ac
          43437 => x"80", -- $0a9ad
          43438 => x"80", -- $0a9ae
          43439 => x"80", -- $0a9af
          43440 => x"80", -- $0a9b0
          43441 => x"80", -- $0a9b1
          43442 => x"80", -- $0a9b2
          43443 => x"80", -- $0a9b3
          43444 => x"80", -- $0a9b4
          43445 => x"80", -- $0a9b5
          43446 => x"80", -- $0a9b6
          43447 => x"80", -- $0a9b7
          43448 => x"80", -- $0a9b8
          43449 => x"80", -- $0a9b9
          43450 => x"80", -- $0a9ba
          43451 => x"80", -- $0a9bb
          43452 => x"80", -- $0a9bc
          43453 => x"80", -- $0a9bd
          43454 => x"80", -- $0a9be
          43455 => x"80", -- $0a9bf
          43456 => x"80", -- $0a9c0
          43457 => x"80", -- $0a9c1
          43458 => x"80", -- $0a9c2
          43459 => x"80", -- $0a9c3
          43460 => x"80", -- $0a9c4
          43461 => x"80", -- $0a9c5
          43462 => x"80", -- $0a9c6
          43463 => x"80", -- $0a9c7
          43464 => x"80", -- $0a9c8
          43465 => x"80", -- $0a9c9
          43466 => x"80", -- $0a9ca
          43467 => x"80", -- $0a9cb
          43468 => x"80", -- $0a9cc
          43469 => x"80", -- $0a9cd
          43470 => x"80", -- $0a9ce
          43471 => x"80", -- $0a9cf
          43472 => x"80", -- $0a9d0
          43473 => x"80", -- $0a9d1
          43474 => x"80", -- $0a9d2
          43475 => x"80", -- $0a9d3
          43476 => x"80", -- $0a9d4
          43477 => x"80", -- $0a9d5
          43478 => x"80", -- $0a9d6
          43479 => x"80", -- $0a9d7
          43480 => x"80", -- $0a9d8
          43481 => x"80", -- $0a9d9
          43482 => x"80", -- $0a9da
          43483 => x"80", -- $0a9db
          43484 => x"80", -- $0a9dc
          43485 => x"80", -- $0a9dd
          43486 => x"7f", -- $0a9de
          43487 => x"7f", -- $0a9df
          43488 => x"7f", -- $0a9e0
          43489 => x"7f", -- $0a9e1
          43490 => x"7f", -- $0a9e2
          43491 => x"7f", -- $0a9e3
          43492 => x"7f", -- $0a9e4
          43493 => x"7f", -- $0a9e5
          43494 => x"7f", -- $0a9e6
          43495 => x"7f", -- $0a9e7
          43496 => x"80", -- $0a9e8
          43497 => x"80", -- $0a9e9
          43498 => x"80", -- $0a9ea
          43499 => x"80", -- $0a9eb
          43500 => x"80", -- $0a9ec
          43501 => x"80", -- $0a9ed
          43502 => x"80", -- $0a9ee
          43503 => x"80", -- $0a9ef
          43504 => x"80", -- $0a9f0
          43505 => x"80", -- $0a9f1
          43506 => x"80", -- $0a9f2
          43507 => x"80", -- $0a9f3
          43508 => x"80", -- $0a9f4
          43509 => x"80", -- $0a9f5
          43510 => x"80", -- $0a9f6
          43511 => x"80", -- $0a9f7
          43512 => x"80", -- $0a9f8
          43513 => x"80", -- $0a9f9
          43514 => x"7f", -- $0a9fa
          43515 => x"7f", -- $0a9fb
          43516 => x"7f", -- $0a9fc
          43517 => x"7f", -- $0a9fd
          43518 => x"7f", -- $0a9fe
          43519 => x"7f", -- $0a9ff
          43520 => x"7f", -- $0aa00
          43521 => x"7f", -- $0aa01
          43522 => x"7f", -- $0aa02
          43523 => x"7f", -- $0aa03
          43524 => x"80", -- $0aa04
          43525 => x"80", -- $0aa05
          43526 => x"80", -- $0aa06
          43527 => x"80", -- $0aa07
          43528 => x"80", -- $0aa08
          43529 => x"80", -- $0aa09
          43530 => x"80", -- $0aa0a
          43531 => x"80", -- $0aa0b
          43532 => x"80", -- $0aa0c
          43533 => x"80", -- $0aa0d
          43534 => x"80", -- $0aa0e
          43535 => x"80", -- $0aa0f
          43536 => x"80", -- $0aa10
          43537 => x"80", -- $0aa11
          43538 => x"80", -- $0aa12
          43539 => x"80", -- $0aa13
          43540 => x"80", -- $0aa14
          43541 => x"80", -- $0aa15
          43542 => x"7f", -- $0aa16
          43543 => x"7f", -- $0aa17
          43544 => x"7f", -- $0aa18
          43545 => x"7f", -- $0aa19
          43546 => x"7f", -- $0aa1a
          43547 => x"7f", -- $0aa1b
          43548 => x"80", -- $0aa1c
          43549 => x"80", -- $0aa1d
          43550 => x"80", -- $0aa1e
          43551 => x"80", -- $0aa1f
          43552 => x"80", -- $0aa20
          43553 => x"80", -- $0aa21
          43554 => x"80", -- $0aa22
          43555 => x"80", -- $0aa23
          43556 => x"80", -- $0aa24
          43557 => x"80", -- $0aa25
          43558 => x"80", -- $0aa26
          43559 => x"80", -- $0aa27
          43560 => x"80", -- $0aa28
          43561 => x"80", -- $0aa29
          43562 => x"80", -- $0aa2a
          43563 => x"80", -- $0aa2b
          43564 => x"80", -- $0aa2c
          43565 => x"80", -- $0aa2d
          43566 => x"80", -- $0aa2e
          43567 => x"7f", -- $0aa2f
          43568 => x"7f", -- $0aa30
          43569 => x"7f", -- $0aa31
          43570 => x"7f", -- $0aa32
          43571 => x"7f", -- $0aa33
          43572 => x"7f", -- $0aa34
          43573 => x"7f", -- $0aa35
          43574 => x"7f", -- $0aa36
          43575 => x"80", -- $0aa37
          43576 => x"80", -- $0aa38
          43577 => x"80", -- $0aa39
          43578 => x"80", -- $0aa3a
          43579 => x"80", -- $0aa3b
          43580 => x"80", -- $0aa3c
          43581 => x"80", -- $0aa3d
          43582 => x"80", -- $0aa3e
          43583 => x"80", -- $0aa3f
          43584 => x"80", -- $0aa40
          43585 => x"80", -- $0aa41
          43586 => x"80", -- $0aa42
          43587 => x"80", -- $0aa43
          43588 => x"80", -- $0aa44
          43589 => x"80", -- $0aa45
          43590 => x"80", -- $0aa46
          43591 => x"7f", -- $0aa47
          43592 => x"7f", -- $0aa48
          43593 => x"7f", -- $0aa49
          43594 => x"7f", -- $0aa4a
          43595 => x"7f", -- $0aa4b
          43596 => x"7f", -- $0aa4c
          43597 => x"7f", -- $0aa4d
          43598 => x"7f", -- $0aa4e
          43599 => x"7f", -- $0aa4f
          43600 => x"7f", -- $0aa50
          43601 => x"7f", -- $0aa51
          43602 => x"7f", -- $0aa52
          43603 => x"7f", -- $0aa53
          43604 => x"7f", -- $0aa54
          43605 => x"7f", -- $0aa55
          43606 => x"7f", -- $0aa56
          43607 => x"80", -- $0aa57
          43608 => x"80", -- $0aa58
          43609 => x"80", -- $0aa59
          43610 => x"80", -- $0aa5a
          43611 => x"80", -- $0aa5b
          43612 => x"80", -- $0aa5c
          43613 => x"80", -- $0aa5d
          43614 => x"7f", -- $0aa5e
          43615 => x"7f", -- $0aa5f
          43616 => x"7f", -- $0aa60
          43617 => x"7f", -- $0aa61
          43618 => x"7f", -- $0aa62
          43619 => x"7f", -- $0aa63
          43620 => x"7f", -- $0aa64
          43621 => x"7f", -- $0aa65
          43622 => x"7f", -- $0aa66
          43623 => x"7f", -- $0aa67
          43624 => x"7f", -- $0aa68
          43625 => x"7f", -- $0aa69
          43626 => x"7f", -- $0aa6a
          43627 => x"7f", -- $0aa6b
          43628 => x"7f", -- $0aa6c
          43629 => x"7f", -- $0aa6d
          43630 => x"7f", -- $0aa6e
          43631 => x"7f", -- $0aa6f
          43632 => x"7f", -- $0aa70
          43633 => x"7f", -- $0aa71
          43634 => x"7f", -- $0aa72
          43635 => x"7f", -- $0aa73
          43636 => x"7f", -- $0aa74
          43637 => x"7f", -- $0aa75
          43638 => x"7f", -- $0aa76
          43639 => x"7f", -- $0aa77
          43640 => x"7f", -- $0aa78
          43641 => x"7f", -- $0aa79
          43642 => x"7f", -- $0aa7a
          43643 => x"7e", -- $0aa7b
          43644 => x"7e", -- $0aa7c
          43645 => x"7e", -- $0aa7d
          43646 => x"7e", -- $0aa7e
          43647 => x"7e", -- $0aa7f
          43648 => x"7e", -- $0aa80
          43649 => x"7e", -- $0aa81
          43650 => x"7e", -- $0aa82
          43651 => x"7e", -- $0aa83
          43652 => x"7f", -- $0aa84
          43653 => x"7f", -- $0aa85
          43654 => x"7f", -- $0aa86
          43655 => x"7f", -- $0aa87
          43656 => x"7f", -- $0aa88
          43657 => x"7f", -- $0aa89
          43658 => x"7f", -- $0aa8a
          43659 => x"7f", -- $0aa8b
          43660 => x"7f", -- $0aa8c
          43661 => x"7f", -- $0aa8d
          43662 => x"7f", -- $0aa8e
          43663 => x"7f", -- $0aa8f
          43664 => x"7f", -- $0aa90
          43665 => x"7f", -- $0aa91
          43666 => x"7f", -- $0aa92
          43667 => x"7e", -- $0aa93
          43668 => x"7e", -- $0aa94
          43669 => x"7e", -- $0aa95
          43670 => x"7e", -- $0aa96
          43671 => x"7e", -- $0aa97
          43672 => x"7e", -- $0aa98
          43673 => x"7f", -- $0aa99
          43674 => x"7f", -- $0aa9a
          43675 => x"7f", -- $0aa9b
          43676 => x"7f", -- $0aa9c
          43677 => x"7f", -- $0aa9d
          43678 => x"7f", -- $0aa9e
          43679 => x"7f", -- $0aa9f
          43680 => x"7f", -- $0aaa0
          43681 => x"80", -- $0aaa1
          43682 => x"80", -- $0aaa2
          43683 => x"80", -- $0aaa3
          43684 => x"80", -- $0aaa4
          43685 => x"80", -- $0aaa5
          43686 => x"80", -- $0aaa6
          43687 => x"80", -- $0aaa7
          43688 => x"80", -- $0aaa8
          43689 => x"7f", -- $0aaa9
          43690 => x"7f", -- $0aaaa
          43691 => x"7f", -- $0aaab
          43692 => x"7f", -- $0aaac
          43693 => x"7f", -- $0aaad
          43694 => x"7f", -- $0aaae
          43695 => x"7f", -- $0aaaf
          43696 => x"7f", -- $0aab0
          43697 => x"7f", -- $0aab1
          43698 => x"7f", -- $0aab2
          43699 => x"7f", -- $0aab3
          43700 => x"7f", -- $0aab4
          43701 => x"80", -- $0aab5
          43702 => x"80", -- $0aab6
          43703 => x"80", -- $0aab7
          43704 => x"80", -- $0aab8
          43705 => x"80", -- $0aab9
          43706 => x"80", -- $0aaba
          43707 => x"80", -- $0aabb
          43708 => x"80", -- $0aabc
          43709 => x"80", -- $0aabd
          43710 => x"80", -- $0aabe
          43711 => x"80", -- $0aabf
          43712 => x"80", -- $0aac0
          43713 => x"80", -- $0aac1
          43714 => x"80", -- $0aac2
          43715 => x"80", -- $0aac3
          43716 => x"80", -- $0aac4
          43717 => x"80", -- $0aac5
          43718 => x"80", -- $0aac6
          43719 => x"80", -- $0aac7
          43720 => x"80", -- $0aac8
          43721 => x"80", -- $0aac9
          43722 => x"80", -- $0aaca
          43723 => x"80", -- $0aacb
          43724 => x"7f", -- $0aacc
          43725 => x"7f", -- $0aacd
          43726 => x"7f", -- $0aace
          43727 => x"7f", -- $0aacf
          43728 => x"7f", -- $0aad0
          43729 => x"80", -- $0aad1
          43730 => x"80", -- $0aad2
          43731 => x"80", -- $0aad3
          43732 => x"80", -- $0aad4
          43733 => x"80", -- $0aad5
          43734 => x"80", -- $0aad6
          43735 => x"80", -- $0aad7
          43736 => x"80", -- $0aad8
          43737 => x"80", -- $0aad9
          43738 => x"80", -- $0aada
          43739 => x"80", -- $0aadb
          43740 => x"80", -- $0aadc
          43741 => x"80", -- $0aadd
          43742 => x"80", -- $0aade
          43743 => x"80", -- $0aadf
          43744 => x"80", -- $0aae0
          43745 => x"80", -- $0aae1
          43746 => x"80", -- $0aae2
          43747 => x"80", -- $0aae3
          43748 => x"80", -- $0aae4
          43749 => x"80", -- $0aae5
          43750 => x"80", -- $0aae6
          43751 => x"80", -- $0aae7
          43752 => x"80", -- $0aae8
          43753 => x"80", -- $0aae9
          43754 => x"80", -- $0aaea
          43755 => x"80", -- $0aaeb
          43756 => x"80", -- $0aaec
          43757 => x"80", -- $0aaed
          43758 => x"80", -- $0aaee
          43759 => x"80", -- $0aaef
          43760 => x"80", -- $0aaf0
          43761 => x"80", -- $0aaf1
          43762 => x"80", -- $0aaf2
          43763 => x"80", -- $0aaf3
          43764 => x"80", -- $0aaf4
          43765 => x"80", -- $0aaf5
          43766 => x"80", -- $0aaf6
          43767 => x"80", -- $0aaf7
          43768 => x"80", -- $0aaf8
          43769 => x"80", -- $0aaf9
          43770 => x"80", -- $0aafa
          43771 => x"80", -- $0aafb
          43772 => x"80", -- $0aafc
          43773 => x"80", -- $0aafd
          43774 => x"80", -- $0aafe
          43775 => x"80", -- $0aaff
          43776 => x"80", -- $0ab00
          43777 => x"80", -- $0ab01
          43778 => x"80", -- $0ab02
          43779 => x"80", -- $0ab03
          43780 => x"80", -- $0ab04
          43781 => x"80", -- $0ab05
          43782 => x"80", -- $0ab06
          43783 => x"80", -- $0ab07
          43784 => x"80", -- $0ab08
          43785 => x"80", -- $0ab09
          43786 => x"80", -- $0ab0a
          43787 => x"80", -- $0ab0b
          43788 => x"80", -- $0ab0c
          43789 => x"80", -- $0ab0d
          43790 => x"80", -- $0ab0e
          43791 => x"80", -- $0ab0f
          43792 => x"80", -- $0ab10
          43793 => x"80", -- $0ab11
          43794 => x"80", -- $0ab12
          43795 => x"80", -- $0ab13
          43796 => x"80", -- $0ab14
          43797 => x"80", -- $0ab15
          43798 => x"80", -- $0ab16
          43799 => x"80", -- $0ab17
          43800 => x"80", -- $0ab18
          43801 => x"80", -- $0ab19
          43802 => x"80", -- $0ab1a
          43803 => x"80", -- $0ab1b
          43804 => x"80", -- $0ab1c
          43805 => x"80", -- $0ab1d
          43806 => x"80", -- $0ab1e
          43807 => x"80", -- $0ab1f
          43808 => x"80", -- $0ab20
          43809 => x"7f", -- $0ab21
          43810 => x"80", -- $0ab22
          43811 => x"7f", -- $0ab23
          43812 => x"7f", -- $0ab24
          43813 => x"80", -- $0ab25
          43814 => x"80", -- $0ab26
          43815 => x"80", -- $0ab27
          43816 => x"80", -- $0ab28
          43817 => x"80", -- $0ab29
          43818 => x"80", -- $0ab2a
          43819 => x"80", -- $0ab2b
          43820 => x"80", -- $0ab2c
          43821 => x"80", -- $0ab2d
          43822 => x"80", -- $0ab2e
          43823 => x"80", -- $0ab2f
          43824 => x"80", -- $0ab30
          43825 => x"80", -- $0ab31
          43826 => x"80", -- $0ab32
          43827 => x"80", -- $0ab33
          43828 => x"80", -- $0ab34
          43829 => x"80", -- $0ab35
          43830 => x"80", -- $0ab36
          43831 => x"80", -- $0ab37
          43832 => x"80", -- $0ab38
          43833 => x"80", -- $0ab39
          43834 => x"7f", -- $0ab3a
          43835 => x"7f", -- $0ab3b
          43836 => x"7f", -- $0ab3c
          43837 => x"7f", -- $0ab3d
          43838 => x"7f", -- $0ab3e
          43839 => x"7f", -- $0ab3f
          43840 => x"80", -- $0ab40
          43841 => x"80", -- $0ab41
          43842 => x"80", -- $0ab42
          43843 => x"80", -- $0ab43
          43844 => x"80", -- $0ab44
          43845 => x"81", -- $0ab45
          43846 => x"81", -- $0ab46
          43847 => x"80", -- $0ab47
          43848 => x"80", -- $0ab48
          43849 => x"81", -- $0ab49
          43850 => x"80", -- $0ab4a
          43851 => x"80", -- $0ab4b
          43852 => x"80", -- $0ab4c
          43853 => x"80", -- $0ab4d
          43854 => x"80", -- $0ab4e
          43855 => x"7f", -- $0ab4f
          43856 => x"80", -- $0ab50
          43857 => x"7f", -- $0ab51
          43858 => x"7e", -- $0ab52
          43859 => x"7f", -- $0ab53
          43860 => x"7e", -- $0ab54
          43861 => x"7e", -- $0ab55
          43862 => x"7e", -- $0ab56
          43863 => x"7e", -- $0ab57
          43864 => x"7f", -- $0ab58
          43865 => x"7e", -- $0ab59
          43866 => x"7d", -- $0ab5a
          43867 => x"7e", -- $0ab5b
          43868 => x"7e", -- $0ab5c
          43869 => x"7e", -- $0ab5d
          43870 => x"7f", -- $0ab5e
          43871 => x"80", -- $0ab5f
          43872 => x"80", -- $0ab60
          43873 => x"80", -- $0ab61
          43874 => x"80", -- $0ab62
          43875 => x"80", -- $0ab63
          43876 => x"80", -- $0ab64
          43877 => x"80", -- $0ab65
          43878 => x"80", -- $0ab66
          43879 => x"80", -- $0ab67
          43880 => x"7f", -- $0ab68
          43881 => x"7e", -- $0ab69
          43882 => x"7e", -- $0ab6a
          43883 => x"7e", -- $0ab6b
          43884 => x"7e", -- $0ab6c
          43885 => x"7e", -- $0ab6d
          43886 => x"7f", -- $0ab6e
          43887 => x"80", -- $0ab6f
          43888 => x"80", -- $0ab70
          43889 => x"81", -- $0ab71
          43890 => x"83", -- $0ab72
          43891 => x"85", -- $0ab73
          43892 => x"87", -- $0ab74
          43893 => x"89", -- $0ab75
          43894 => x"8a", -- $0ab76
          43895 => x"8b", -- $0ab77
          43896 => x"8c", -- $0ab78
          43897 => x"8d", -- $0ab79
          43898 => x"8d", -- $0ab7a
          43899 => x"8c", -- $0ab7b
          43900 => x"8b", -- $0ab7c
          43901 => x"89", -- $0ab7d
          43902 => x"88", -- $0ab7e
          43903 => x"86", -- $0ab7f
          43904 => x"85", -- $0ab80
          43905 => x"83", -- $0ab81
          43906 => x"82", -- $0ab82
          43907 => x"82", -- $0ab83
          43908 => x"81", -- $0ab84
          43909 => x"81", -- $0ab85
          43910 => x"82", -- $0ab86
          43911 => x"83", -- $0ab87
          43912 => x"84", -- $0ab88
          43913 => x"84", -- $0ab89
          43914 => x"85", -- $0ab8a
          43915 => x"84", -- $0ab8b
          43916 => x"85", -- $0ab8c
          43917 => x"85", -- $0ab8d
          43918 => x"84", -- $0ab8e
          43919 => x"84", -- $0ab8f
          43920 => x"83", -- $0ab90
          43921 => x"83", -- $0ab91
          43922 => x"82", -- $0ab92
          43923 => x"82", -- $0ab93
          43924 => x"82", -- $0ab94
          43925 => x"82", -- $0ab95
          43926 => x"81", -- $0ab96
          43927 => x"81", -- $0ab97
          43928 => x"81", -- $0ab98
          43929 => x"80", -- $0ab99
          43930 => x"80", -- $0ab9a
          43931 => x"80", -- $0ab9b
          43932 => x"7f", -- $0ab9c
          43933 => x"7e", -- $0ab9d
          43934 => x"7d", -- $0ab9e
          43935 => x"7c", -- $0ab9f
          43936 => x"7b", -- $0aba0
          43937 => x"7a", -- $0aba1
          43938 => x"7a", -- $0aba2
          43939 => x"79", -- $0aba3
          43940 => x"78", -- $0aba4
          43941 => x"79", -- $0aba5
          43942 => x"79", -- $0aba6
          43943 => x"79", -- $0aba7
          43944 => x"79", -- $0aba8
          43945 => x"7a", -- $0aba9
          43946 => x"7b", -- $0abaa
          43947 => x"7c", -- $0abab
          43948 => x"7c", -- $0abac
          43949 => x"7d", -- $0abad
          43950 => x"7d", -- $0abae
          43951 => x"7e", -- $0abaf
          43952 => x"7d", -- $0abb0
          43953 => x"7c", -- $0abb1
          43954 => x"7c", -- $0abb2
          43955 => x"7b", -- $0abb3
          43956 => x"7a", -- $0abb4
          43957 => x"79", -- $0abb5
          43958 => x"78", -- $0abb6
          43959 => x"78", -- $0abb7
          43960 => x"78", -- $0abb8
          43961 => x"77", -- $0abb9
          43962 => x"77", -- $0abba
          43963 => x"78", -- $0abbb
          43964 => x"78", -- $0abbc
          43965 => x"78", -- $0abbd
          43966 => x"79", -- $0abbe
          43967 => x"7a", -- $0abbf
          43968 => x"7a", -- $0abc0
          43969 => x"7b", -- $0abc1
          43970 => x"7c", -- $0abc2
          43971 => x"7d", -- $0abc3
          43972 => x"7e", -- $0abc4
          43973 => x"7f", -- $0abc5
          43974 => x"80", -- $0abc6
          43975 => x"80", -- $0abc7
          43976 => x"81", -- $0abc8
          43977 => x"83", -- $0abc9
          43978 => x"84", -- $0abca
          43979 => x"85", -- $0abcb
          43980 => x"86", -- $0abcc
          43981 => x"87", -- $0abcd
          43982 => x"88", -- $0abce
          43983 => x"89", -- $0abcf
          43984 => x"89", -- $0abd0
          43985 => x"89", -- $0abd1
          43986 => x"89", -- $0abd2
          43987 => x"88", -- $0abd3
          43988 => x"88", -- $0abd4
          43989 => x"88", -- $0abd5
          43990 => x"88", -- $0abd6
          43991 => x"88", -- $0abd7
          43992 => x"88", -- $0abd8
          43993 => x"88", -- $0abd9
          43994 => x"88", -- $0abda
          43995 => x"88", -- $0abdb
          43996 => x"88", -- $0abdc
          43997 => x"89", -- $0abdd
          43998 => x"8a", -- $0abde
          43999 => x"8a", -- $0abdf
          44000 => x"8a", -- $0abe0
          44001 => x"8a", -- $0abe1
          44002 => x"89", -- $0abe2
          44003 => x"89", -- $0abe3
          44004 => x"89", -- $0abe4
          44005 => x"88", -- $0abe5
          44006 => x"87", -- $0abe6
          44007 => x"86", -- $0abe7
          44008 => x"86", -- $0abe8
          44009 => x"85", -- $0abe9
          44010 => x"84", -- $0abea
          44011 => x"84", -- $0abeb
          44012 => x"84", -- $0abec
          44013 => x"83", -- $0abed
          44014 => x"83", -- $0abee
          44015 => x"83", -- $0abef
          44016 => x"83", -- $0abf0
          44017 => x"83", -- $0abf1
          44018 => x"82", -- $0abf2
          44019 => x"82", -- $0abf3
          44020 => x"82", -- $0abf4
          44021 => x"81", -- $0abf5
          44022 => x"80", -- $0abf6
          44023 => x"80", -- $0abf7
          44024 => x"80", -- $0abf8
          44025 => x"80", -- $0abf9
          44026 => x"80", -- $0abfa
          44027 => x"80", -- $0abfb
          44028 => x"80", -- $0abfc
          44029 => x"81", -- $0abfd
          44030 => x"82", -- $0abfe
          44031 => x"82", -- $0abff
          44032 => x"82", -- $0ac00
          44033 => x"83", -- $0ac01
          44034 => x"83", -- $0ac02
          44035 => x"83", -- $0ac03
          44036 => x"82", -- $0ac04
          44037 => x"82", -- $0ac05
          44038 => x"81", -- $0ac06
          44039 => x"80", -- $0ac07
          44040 => x"80", -- $0ac08
          44041 => x"7f", -- $0ac09
          44042 => x"7e", -- $0ac0a
          44043 => x"7d", -- $0ac0b
          44044 => x"7c", -- $0ac0c
          44045 => x"7b", -- $0ac0d
          44046 => x"7a", -- $0ac0e
          44047 => x"7a", -- $0ac0f
          44048 => x"7a", -- $0ac10
          44049 => x"7a", -- $0ac11
          44050 => x"7a", -- $0ac12
          44051 => x"7a", -- $0ac13
          44052 => x"7b", -- $0ac14
          44053 => x"7b", -- $0ac15
          44054 => x"7b", -- $0ac16
          44055 => x"7c", -- $0ac17
          44056 => x"7c", -- $0ac18
          44057 => x"7c", -- $0ac19
          44058 => x"7c", -- $0ac1a
          44059 => x"7c", -- $0ac1b
          44060 => x"7c", -- $0ac1c
          44061 => x"7c", -- $0ac1d
          44062 => x"7c", -- $0ac1e
          44063 => x"7d", -- $0ac1f
          44064 => x"7d", -- $0ac20
          44065 => x"7d", -- $0ac21
          44066 => x"7d", -- $0ac22
          44067 => x"7d", -- $0ac23
          44068 => x"7e", -- $0ac24
          44069 => x"7e", -- $0ac25
          44070 => x"7e", -- $0ac26
          44071 => x"7e", -- $0ac27
          44072 => x"7e", -- $0ac28
          44073 => x"7e", -- $0ac29
          44074 => x"7f", -- $0ac2a
          44075 => x"7f", -- $0ac2b
          44076 => x"7f", -- $0ac2c
          44077 => x"80", -- $0ac2d
          44078 => x"80", -- $0ac2e
          44079 => x"80", -- $0ac2f
          44080 => x"80", -- $0ac30
          44081 => x"81", -- $0ac31
          44082 => x"81", -- $0ac32
          44083 => x"81", -- $0ac33
          44084 => x"82", -- $0ac34
          44085 => x"82", -- $0ac35
          44086 => x"83", -- $0ac36
          44087 => x"83", -- $0ac37
          44088 => x"83", -- $0ac38
          44089 => x"83", -- $0ac39
          44090 => x"83", -- $0ac3a
          44091 => x"83", -- $0ac3b
          44092 => x"83", -- $0ac3c
          44093 => x"82", -- $0ac3d
          44094 => x"82", -- $0ac3e
          44095 => x"81", -- $0ac3f
          44096 => x"81", -- $0ac40
          44097 => x"81", -- $0ac41
          44098 => x"81", -- $0ac42
          44099 => x"81", -- $0ac43
          44100 => x"81", -- $0ac44
          44101 => x"81", -- $0ac45
          44102 => x"81", -- $0ac46
          44103 => x"82", -- $0ac47
          44104 => x"82", -- $0ac48
          44105 => x"82", -- $0ac49
          44106 => x"83", -- $0ac4a
          44107 => x"83", -- $0ac4b
          44108 => x"83", -- $0ac4c
          44109 => x"84", -- $0ac4d
          44110 => x"00", -- $0ac4e
          44111 => x"00", -- $0ac4f
          44112 => x"00", -- $0ac50
          44113 => x"00", -- $0ac51
          44114 => x"00", -- $0ac52
          44115 => x"00", -- $0ac53
          44116 => x"00", -- $0ac54
          44117 => x"00", -- $0ac55
          44118 => x"00", -- $0ac56
          44119 => x"00", -- $0ac57
          44120 => x"00", -- $0ac58
          44121 => x"00", -- $0ac59
          44122 => x"00", -- $0ac5a
          44123 => x"00", -- $0ac5b
          44124 => x"00", -- $0ac5c
          44125 => x"00", -- $0ac5d
          44126 => x"00", -- $0ac5e
          44127 => x"00", -- $0ac5f
          44128 => x"00", -- $0ac60
          44129 => x"00", -- $0ac61
          44130 => x"00", -- $0ac62
          44131 => x"00", -- $0ac63
          44132 => x"00", -- $0ac64
          44133 => x"00", -- $0ac65
          44134 => x"00", -- $0ac66
          44135 => x"00", -- $0ac67
          44136 => x"00", -- $0ac68
          44137 => x"00", -- $0ac69
          44138 => x"00", -- $0ac6a
          44139 => x"00", -- $0ac6b
          44140 => x"00", -- $0ac6c
          44141 => x"00", -- $0ac6d
          44142 => x"00", -- $0ac6e
          44143 => x"00", -- $0ac6f
          44144 => x"00", -- $0ac70
          44145 => x"00", -- $0ac71
          44146 => x"00", -- $0ac72
          44147 => x"00", -- $0ac73
          44148 => x"00", -- $0ac74
          44149 => x"00", -- $0ac75
          44150 => x"00", -- $0ac76
          44151 => x"00", -- $0ac77
          44152 => x"00", -- $0ac78
          44153 => x"00", -- $0ac79
          44154 => x"00", -- $0ac7a
          44155 => x"00", -- $0ac7b
          44156 => x"00", -- $0ac7c
          44157 => x"00", -- $0ac7d
          44158 => x"00", -- $0ac7e
          44159 => x"00", -- $0ac7f
          44160 => x"00", -- $0ac80
          44161 => x"00", -- $0ac81
          44162 => x"00", -- $0ac82
          44163 => x"00", -- $0ac83
          44164 => x"00", -- $0ac84
          44165 => x"00", -- $0ac85
          44166 => x"00", -- $0ac86
          44167 => x"00", -- $0ac87
          44168 => x"00", -- $0ac88
          44169 => x"00", -- $0ac89
          44170 => x"00", -- $0ac8a
          44171 => x"00", -- $0ac8b
          44172 => x"00", -- $0ac8c
          44173 => x"00", -- $0ac8d
          44174 => x"00", -- $0ac8e
          44175 => x"00", -- $0ac8f
          44176 => x"00", -- $0ac90
          44177 => x"00", -- $0ac91
          44178 => x"00", -- $0ac92
          44179 => x"00", -- $0ac93
          44180 => x"00", -- $0ac94
          44181 => x"00", -- $0ac95
          44182 => x"00", -- $0ac96
          44183 => x"00", -- $0ac97
          44184 => x"00", -- $0ac98
          44185 => x"00", -- $0ac99
          44186 => x"00", -- $0ac9a
          44187 => x"00", -- $0ac9b
          44188 => x"00", -- $0ac9c
          44189 => x"00", -- $0ac9d
          44190 => x"00", -- $0ac9e
          44191 => x"00", -- $0ac9f
          44192 => x"00", -- $0aca0
          44193 => x"00", -- $0aca1
          44194 => x"00", -- $0aca2
          44195 => x"00", -- $0aca3
          44196 => x"00", -- $0aca4
          44197 => x"00", -- $0aca5
          44198 => x"00", -- $0aca6
          44199 => x"00", -- $0aca7
          44200 => x"00", -- $0aca8
          44201 => x"00", -- $0aca9
          44202 => x"00", -- $0acaa
          44203 => x"00", -- $0acab
          44204 => x"00", -- $0acac
          44205 => x"00", -- $0acad
          44206 => x"00", -- $0acae
          44207 => x"00", -- $0acaf
          44208 => x"00", -- $0acb0
          44209 => x"00", -- $0acb1
          44210 => x"00", -- $0acb2
          44211 => x"00", -- $0acb3
          44212 => x"00", -- $0acb4
          44213 => x"00", -- $0acb5
          44214 => x"00", -- $0acb6
          44215 => x"00", -- $0acb7
          44216 => x"00", -- $0acb8
          44217 => x"00", -- $0acb9
          44218 => x"00", -- $0acba
          44219 => x"00", -- $0acbb
          44220 => x"00", -- $0acbc
          44221 => x"00", -- $0acbd
          44222 => x"00", -- $0acbe
          44223 => x"00", -- $0acbf
          44224 => x"00", -- $0acc0
          44225 => x"00", -- $0acc1
          44226 => x"00", -- $0acc2
          44227 => x"00", -- $0acc3
          44228 => x"00", -- $0acc4
          44229 => x"00", -- $0acc5
          44230 => x"00", -- $0acc6
          44231 => x"00", -- $0acc7
          44232 => x"00", -- $0acc8
          44233 => x"00", -- $0acc9
          44234 => x"00", -- $0acca
          44235 => x"00", -- $0accb
          44236 => x"00", -- $0accc
          44237 => x"00", -- $0accd
          44238 => x"00", -- $0acce
          44239 => x"00", -- $0accf
          44240 => x"00", -- $0acd0
          44241 => x"00", -- $0acd1
          44242 => x"00", -- $0acd2
          44243 => x"00", -- $0acd3
          44244 => x"00", -- $0acd4
          44245 => x"00", -- $0acd5
          44246 => x"00", -- $0acd6
          44247 => x"00", -- $0acd7
          44248 => x"00", -- $0acd8
          44249 => x"00", -- $0acd9
          44250 => x"00", -- $0acda
          44251 => x"00", -- $0acdb
          44252 => x"00", -- $0acdc
          44253 => x"00", -- $0acdd
          44254 => x"00", -- $0acde
          44255 => x"00", -- $0acdf
          44256 => x"00", -- $0ace0
          44257 => x"00", -- $0ace1
          44258 => x"00", -- $0ace2
          44259 => x"00", -- $0ace3
          44260 => x"00", -- $0ace4
          44261 => x"00", -- $0ace5
          44262 => x"00", -- $0ace6
          44263 => x"00", -- $0ace7
          44264 => x"00", -- $0ace8
          44265 => x"00", -- $0ace9
          44266 => x"00", -- $0acea
          44267 => x"00", -- $0aceb
          44268 => x"00", -- $0acec
          44269 => x"00", -- $0aced
          44270 => x"00", -- $0acee
          44271 => x"00", -- $0acef
          44272 => x"00", -- $0acf0
          44273 => x"00", -- $0acf1
          44274 => x"00", -- $0acf2
          44275 => x"00", -- $0acf3
          44276 => x"00", -- $0acf4
          44277 => x"00", -- $0acf5
          44278 => x"00", -- $0acf6
          44279 => x"00", -- $0acf7
          44280 => x"00", -- $0acf8
          44281 => x"00", -- $0acf9
          44282 => x"00", -- $0acfa
          44283 => x"00", -- $0acfb
          44284 => x"00", -- $0acfc
          44285 => x"00", -- $0acfd
          44286 => x"00", -- $0acfe
          44287 => x"00", -- $0acff
          44288 => x"00", -- $0ad00
          44289 => x"00", -- $0ad01
          44290 => x"00", -- $0ad02
          44291 => x"00", -- $0ad03
          44292 => x"00", -- $0ad04
          44293 => x"00", -- $0ad05
          44294 => x"00", -- $0ad06
          44295 => x"00", -- $0ad07
          44296 => x"00", -- $0ad08
          44297 => x"00", -- $0ad09
          44298 => x"00", -- $0ad0a
          44299 => x"00", -- $0ad0b
          44300 => x"00", -- $0ad0c
          44301 => x"00", -- $0ad0d
          44302 => x"00", -- $0ad0e
          44303 => x"00", -- $0ad0f
          44304 => x"00", -- $0ad10
          44305 => x"00", -- $0ad11
          44306 => x"00", -- $0ad12
          44307 => x"00", -- $0ad13
          44308 => x"00", -- $0ad14
          44309 => x"00", -- $0ad15
          44310 => x"00", -- $0ad16
          44311 => x"00", -- $0ad17
          44312 => x"00", -- $0ad18
          44313 => x"00", -- $0ad19
          44314 => x"00", -- $0ad1a
          44315 => x"00", -- $0ad1b
          44316 => x"00", -- $0ad1c
          44317 => x"00", -- $0ad1d
          44318 => x"00", -- $0ad1e
          44319 => x"00", -- $0ad1f
          44320 => x"00", -- $0ad20
          44321 => x"00", -- $0ad21
          44322 => x"00", -- $0ad22
          44323 => x"00", -- $0ad23
          44324 => x"00", -- $0ad24
          44325 => x"00", -- $0ad25
          44326 => x"00", -- $0ad26
          44327 => x"00", -- $0ad27
          44328 => x"00", -- $0ad28
          44329 => x"00", -- $0ad29
          44330 => x"00", -- $0ad2a
          44331 => x"00", -- $0ad2b
          44332 => x"00", -- $0ad2c
          44333 => x"00", -- $0ad2d
          44334 => x"00", -- $0ad2e
          44335 => x"00", -- $0ad2f
          44336 => x"00", -- $0ad30
          44337 => x"00", -- $0ad31
          44338 => x"00", -- $0ad32
          44339 => x"00", -- $0ad33
          44340 => x"00", -- $0ad34
          44341 => x"00", -- $0ad35
          44342 => x"00", -- $0ad36
          44343 => x"00", -- $0ad37
          44344 => x"00", -- $0ad38
          44345 => x"00", -- $0ad39
          44346 => x"00", -- $0ad3a
          44347 => x"00", -- $0ad3b
          44348 => x"00", -- $0ad3c
          44349 => x"00", -- $0ad3d
          44350 => x"00", -- $0ad3e
          44351 => x"00", -- $0ad3f
          44352 => x"00", -- $0ad40
          44353 => x"00", -- $0ad41
          44354 => x"00", -- $0ad42
          44355 => x"00", -- $0ad43
          44356 => x"00", -- $0ad44
          44357 => x"00", -- $0ad45
          44358 => x"00", -- $0ad46
          44359 => x"00", -- $0ad47
          44360 => x"00", -- $0ad48
          44361 => x"00", -- $0ad49
          44362 => x"00", -- $0ad4a
          44363 => x"00", -- $0ad4b
          44364 => x"00", -- $0ad4c
          44365 => x"00", -- $0ad4d
          44366 => x"00", -- $0ad4e
          44367 => x"00", -- $0ad4f
          44368 => x"00", -- $0ad50
          44369 => x"00", -- $0ad51
          44370 => x"00", -- $0ad52
          44371 => x"00", -- $0ad53
          44372 => x"00", -- $0ad54
          44373 => x"00", -- $0ad55
          44374 => x"00", -- $0ad56
          44375 => x"00", -- $0ad57
          44376 => x"00", -- $0ad58
          44377 => x"00", -- $0ad59
          44378 => x"00", -- $0ad5a
          44379 => x"00", -- $0ad5b
          44380 => x"00", -- $0ad5c
          44381 => x"00", -- $0ad5d
          44382 => x"00", -- $0ad5e
          44383 => x"00", -- $0ad5f
          44384 => x"00", -- $0ad60
          44385 => x"00", -- $0ad61
          44386 => x"00", -- $0ad62
          44387 => x"00", -- $0ad63
          44388 => x"00", -- $0ad64
          44389 => x"00", -- $0ad65
          44390 => x"00", -- $0ad66
          44391 => x"00", -- $0ad67
          44392 => x"00", -- $0ad68
          44393 => x"00", -- $0ad69
          44394 => x"00", -- $0ad6a
          44395 => x"00", -- $0ad6b
          44396 => x"00", -- $0ad6c
          44397 => x"00", -- $0ad6d
          44398 => x"00", -- $0ad6e
          44399 => x"00", -- $0ad6f
          44400 => x"00", -- $0ad70
          44401 => x"00", -- $0ad71
          44402 => x"00", -- $0ad72
          44403 => x"00", -- $0ad73
          44404 => x"00", -- $0ad74
          44405 => x"00", -- $0ad75
          44406 => x"00", -- $0ad76
          44407 => x"00", -- $0ad77
          44408 => x"00", -- $0ad78
          44409 => x"00", -- $0ad79
          44410 => x"00", -- $0ad7a
          44411 => x"00", -- $0ad7b
          44412 => x"00", -- $0ad7c
          44413 => x"00", -- $0ad7d
          44414 => x"00", -- $0ad7e
          44415 => x"00", -- $0ad7f
          44416 => x"00", -- $0ad80
          44417 => x"00", -- $0ad81
          44418 => x"00", -- $0ad82
          44419 => x"00", -- $0ad83
          44420 => x"00", -- $0ad84
          44421 => x"00", -- $0ad85
          44422 => x"00", -- $0ad86
          44423 => x"00", -- $0ad87
          44424 => x"00", -- $0ad88
          44425 => x"00", -- $0ad89
          44426 => x"00", -- $0ad8a
          44427 => x"00", -- $0ad8b
          44428 => x"00", -- $0ad8c
          44429 => x"00", -- $0ad8d
          44430 => x"00", -- $0ad8e
          44431 => x"00", -- $0ad8f
          44432 => x"00", -- $0ad90
          44433 => x"00", -- $0ad91
          44434 => x"00", -- $0ad92
          44435 => x"00", -- $0ad93
          44436 => x"00", -- $0ad94
          44437 => x"00", -- $0ad95
          44438 => x"00", -- $0ad96
          44439 => x"00", -- $0ad97
          44440 => x"00", -- $0ad98
          44441 => x"00", -- $0ad99
          44442 => x"00", -- $0ad9a
          44443 => x"00", -- $0ad9b
          44444 => x"00", -- $0ad9c
          44445 => x"00", -- $0ad9d
          44446 => x"00", -- $0ad9e
          44447 => x"00", -- $0ad9f
          44448 => x"00", -- $0ada0
          44449 => x"00", -- $0ada1
          44450 => x"00", -- $0ada2
          44451 => x"00", -- $0ada3
          44452 => x"00", -- $0ada4
          44453 => x"00", -- $0ada5
          44454 => x"00", -- $0ada6
          44455 => x"00", -- $0ada7
          44456 => x"00", -- $0ada8
          44457 => x"00", -- $0ada9
          44458 => x"00", -- $0adaa
          44459 => x"00", -- $0adab
          44460 => x"00", -- $0adac
          44461 => x"00", -- $0adad
          44462 => x"00", -- $0adae
          44463 => x"00", -- $0adaf
          44464 => x"00", -- $0adb0
          44465 => x"00", -- $0adb1
          44466 => x"00", -- $0adb2
          44467 => x"00", -- $0adb3
          44468 => x"00", -- $0adb4
          44469 => x"00", -- $0adb5
          44470 => x"00", -- $0adb6
          44471 => x"00", -- $0adb7
          44472 => x"00", -- $0adb8
          44473 => x"00", -- $0adb9
          44474 => x"00", -- $0adba
          44475 => x"00", -- $0adbb
          44476 => x"00", -- $0adbc
          44477 => x"00", -- $0adbd
          44478 => x"00", -- $0adbe
          44479 => x"00", -- $0adbf
          44480 => x"00", -- $0adc0
          44481 => x"00", -- $0adc1
          44482 => x"00", -- $0adc2
          44483 => x"00", -- $0adc3
          44484 => x"00", -- $0adc4
          44485 => x"00", -- $0adc5
          44486 => x"00", -- $0adc6
          44487 => x"00", -- $0adc7
          44488 => x"00", -- $0adc8
          44489 => x"00", -- $0adc9
          44490 => x"00", -- $0adca
          44491 => x"00", -- $0adcb
          44492 => x"00", -- $0adcc
          44493 => x"00", -- $0adcd
          44494 => x"00", -- $0adce
          44495 => x"00", -- $0adcf
          44496 => x"00", -- $0add0
          44497 => x"00", -- $0add1
          44498 => x"00", -- $0add2
          44499 => x"00", -- $0add3
          44500 => x"00", -- $0add4
          44501 => x"00", -- $0add5
          44502 => x"00", -- $0add6
          44503 => x"00", -- $0add7
          44504 => x"00", -- $0add8
          44505 => x"00", -- $0add9
          44506 => x"00", -- $0adda
          44507 => x"00", -- $0addb
          44508 => x"00", -- $0addc
          44509 => x"00", -- $0addd
          44510 => x"00", -- $0adde
          44511 => x"00", -- $0addf
          44512 => x"00", -- $0ade0
          44513 => x"00", -- $0ade1
          44514 => x"00", -- $0ade2
          44515 => x"00", -- $0ade3
          44516 => x"00", -- $0ade4
          44517 => x"00", -- $0ade5
          44518 => x"00", -- $0ade6
          44519 => x"00", -- $0ade7
          44520 => x"00", -- $0ade8
          44521 => x"00", -- $0ade9
          44522 => x"00", -- $0adea
          44523 => x"00", -- $0adeb
          44524 => x"00", -- $0adec
          44525 => x"00", -- $0aded
          44526 => x"00", -- $0adee
          44527 => x"00", -- $0adef
          44528 => x"00", -- $0adf0
          44529 => x"00", -- $0adf1
          44530 => x"00", -- $0adf2
          44531 => x"00", -- $0adf3
          44532 => x"00", -- $0adf4
          44533 => x"00", -- $0adf5
          44534 => x"00", -- $0adf6
          44535 => x"00", -- $0adf7
          44536 => x"00", -- $0adf8
          44537 => x"00", -- $0adf9
          44538 => x"00", -- $0adfa
          44539 => x"00", -- $0adfb
          44540 => x"00", -- $0adfc
          44541 => x"00", -- $0adfd
          44542 => x"00", -- $0adfe
          44543 => x"00", -- $0adff
          44544 => x"00", -- $0ae00
          44545 => x"00", -- $0ae01
          44546 => x"00", -- $0ae02
          44547 => x"00", -- $0ae03
          44548 => x"00", -- $0ae04
          44549 => x"00", -- $0ae05
          44550 => x"00", -- $0ae06
          44551 => x"00", -- $0ae07
          44552 => x"00", -- $0ae08
          44553 => x"00", -- $0ae09
          44554 => x"00", -- $0ae0a
          44555 => x"00", -- $0ae0b
          44556 => x"00", -- $0ae0c
          44557 => x"00", -- $0ae0d
          44558 => x"00", -- $0ae0e
          44559 => x"00", -- $0ae0f
          44560 => x"00", -- $0ae10
          44561 => x"00", -- $0ae11
          44562 => x"00", -- $0ae12
          44563 => x"00", -- $0ae13
          44564 => x"00", -- $0ae14
          44565 => x"00", -- $0ae15
          44566 => x"00", -- $0ae16
          44567 => x"00", -- $0ae17
          44568 => x"00", -- $0ae18
          44569 => x"00", -- $0ae19
          44570 => x"00", -- $0ae1a
          44571 => x"00", -- $0ae1b
          44572 => x"00", -- $0ae1c
          44573 => x"00", -- $0ae1d
          44574 => x"00", -- $0ae1e
          44575 => x"00", -- $0ae1f
          44576 => x"00", -- $0ae20
          44577 => x"00", -- $0ae21
          44578 => x"00", -- $0ae22
          44579 => x"00", -- $0ae23
          44580 => x"00", -- $0ae24
          44581 => x"00", -- $0ae25
          44582 => x"00", -- $0ae26
          44583 => x"00", -- $0ae27
          44584 => x"00", -- $0ae28
          44585 => x"00", -- $0ae29
          44586 => x"00", -- $0ae2a
          44587 => x"00", -- $0ae2b
          44588 => x"00", -- $0ae2c
          44589 => x"00", -- $0ae2d
          44590 => x"00", -- $0ae2e
          44591 => x"00", -- $0ae2f
          44592 => x"00", -- $0ae30
          44593 => x"00", -- $0ae31
          44594 => x"00", -- $0ae32
          44595 => x"00", -- $0ae33
          44596 => x"00", -- $0ae34
          44597 => x"00", -- $0ae35
          44598 => x"00", -- $0ae36
          44599 => x"00", -- $0ae37
          44600 => x"00", -- $0ae38
          44601 => x"00", -- $0ae39
          44602 => x"00", -- $0ae3a
          44603 => x"00", -- $0ae3b
          44604 => x"00", -- $0ae3c
          44605 => x"00", -- $0ae3d
          44606 => x"00", -- $0ae3e
          44607 => x"00", -- $0ae3f
          44608 => x"00", -- $0ae40
          44609 => x"00", -- $0ae41
          44610 => x"00", -- $0ae42
          44611 => x"00", -- $0ae43
          44612 => x"00", -- $0ae44
          44613 => x"00", -- $0ae45
          44614 => x"00", -- $0ae46
          44615 => x"00", -- $0ae47
          44616 => x"00", -- $0ae48
          44617 => x"00", -- $0ae49
          44618 => x"00", -- $0ae4a
          44619 => x"00", -- $0ae4b
          44620 => x"00", -- $0ae4c
          44621 => x"00", -- $0ae4d
          44622 => x"00", -- $0ae4e
          44623 => x"00", -- $0ae4f
          44624 => x"00", -- $0ae50
          44625 => x"00", -- $0ae51
          44626 => x"00", -- $0ae52
          44627 => x"00", -- $0ae53
          44628 => x"00", -- $0ae54
          44629 => x"00", -- $0ae55
          44630 => x"00", -- $0ae56
          44631 => x"00", -- $0ae57
          44632 => x"00", -- $0ae58
          44633 => x"00", -- $0ae59
          44634 => x"00", -- $0ae5a
          44635 => x"00", -- $0ae5b
          44636 => x"00", -- $0ae5c
          44637 => x"00", -- $0ae5d
          44638 => x"00", -- $0ae5e
          44639 => x"00", -- $0ae5f
          44640 => x"00", -- $0ae60
          44641 => x"00", -- $0ae61
          44642 => x"00", -- $0ae62
          44643 => x"00", -- $0ae63
          44644 => x"00", -- $0ae64
          44645 => x"00", -- $0ae65
          44646 => x"00", -- $0ae66
          44647 => x"00", -- $0ae67
          44648 => x"00", -- $0ae68
          44649 => x"00", -- $0ae69
          44650 => x"00", -- $0ae6a
          44651 => x"00", -- $0ae6b
          44652 => x"00", -- $0ae6c
          44653 => x"00", -- $0ae6d
          44654 => x"00", -- $0ae6e
          44655 => x"00", -- $0ae6f
          44656 => x"00", -- $0ae70
          44657 => x"00", -- $0ae71
          44658 => x"00", -- $0ae72
          44659 => x"00", -- $0ae73
          44660 => x"00", -- $0ae74
          44661 => x"00", -- $0ae75
          44662 => x"00", -- $0ae76
          44663 => x"00", -- $0ae77
          44664 => x"00", -- $0ae78
          44665 => x"00", -- $0ae79
          44666 => x"00", -- $0ae7a
          44667 => x"00", -- $0ae7b
          44668 => x"00", -- $0ae7c
          44669 => x"00", -- $0ae7d
          44670 => x"00", -- $0ae7e
          44671 => x"00", -- $0ae7f
          44672 => x"00", -- $0ae80
          44673 => x"00", -- $0ae81
          44674 => x"00", -- $0ae82
          44675 => x"00", -- $0ae83
          44676 => x"00", -- $0ae84
          44677 => x"00", -- $0ae85
          44678 => x"00", -- $0ae86
          44679 => x"00", -- $0ae87
          44680 => x"00", -- $0ae88
          44681 => x"00", -- $0ae89
          44682 => x"00", -- $0ae8a
          44683 => x"00", -- $0ae8b
          44684 => x"00", -- $0ae8c
          44685 => x"00", -- $0ae8d
          44686 => x"00", -- $0ae8e
          44687 => x"00", -- $0ae8f
          44688 => x"00", -- $0ae90
          44689 => x"00", -- $0ae91
          44690 => x"00", -- $0ae92
          44691 => x"00", -- $0ae93
          44692 => x"00", -- $0ae94
          44693 => x"00", -- $0ae95
          44694 => x"00", -- $0ae96
          44695 => x"00", -- $0ae97
          44696 => x"00", -- $0ae98
          44697 => x"00", -- $0ae99
          44698 => x"00", -- $0ae9a
          44699 => x"00", -- $0ae9b
          44700 => x"00", -- $0ae9c
          44701 => x"00", -- $0ae9d
          44702 => x"00", -- $0ae9e
          44703 => x"00", -- $0ae9f
          44704 => x"00", -- $0aea0
          44705 => x"00", -- $0aea1
          44706 => x"00", -- $0aea2
          44707 => x"00", -- $0aea3
          44708 => x"00", -- $0aea4
          44709 => x"00", -- $0aea5
          44710 => x"00", -- $0aea6
          44711 => x"00", -- $0aea7
          44712 => x"00", -- $0aea8
          44713 => x"00", -- $0aea9
          44714 => x"00", -- $0aeaa
          44715 => x"00", -- $0aeab
          44716 => x"00", -- $0aeac
          44717 => x"00", -- $0aead
          44718 => x"00", -- $0aeae
          44719 => x"00", -- $0aeaf
          44720 => x"00", -- $0aeb0
          44721 => x"00", -- $0aeb1
          44722 => x"00", -- $0aeb2
          44723 => x"00", -- $0aeb3
          44724 => x"00", -- $0aeb4
          44725 => x"00", -- $0aeb5
          44726 => x"00", -- $0aeb6
          44727 => x"00", -- $0aeb7
          44728 => x"00", -- $0aeb8
          44729 => x"00", -- $0aeb9
          44730 => x"00", -- $0aeba
          44731 => x"00", -- $0aebb
          44732 => x"00", -- $0aebc
          44733 => x"00", -- $0aebd
          44734 => x"00", -- $0aebe
          44735 => x"00", -- $0aebf
          44736 => x"00", -- $0aec0
          44737 => x"00", -- $0aec1
          44738 => x"00", -- $0aec2
          44739 => x"00", -- $0aec3
          44740 => x"00", -- $0aec4
          44741 => x"00", -- $0aec5
          44742 => x"00", -- $0aec6
          44743 => x"00", -- $0aec7
          44744 => x"00", -- $0aec8
          44745 => x"00", -- $0aec9
          44746 => x"00", -- $0aeca
          44747 => x"00", -- $0aecb
          44748 => x"00", -- $0aecc
          44749 => x"00", -- $0aecd
          44750 => x"00", -- $0aece
          44751 => x"00", -- $0aecf
          44752 => x"00", -- $0aed0
          44753 => x"00", -- $0aed1
          44754 => x"00", -- $0aed2
          44755 => x"00", -- $0aed3
          44756 => x"00", -- $0aed4
          44757 => x"00", -- $0aed5
          44758 => x"00", -- $0aed6
          44759 => x"00", -- $0aed7
          44760 => x"00", -- $0aed8
          44761 => x"00", -- $0aed9
          44762 => x"00", -- $0aeda
          44763 => x"00", -- $0aedb
          44764 => x"00", -- $0aedc
          44765 => x"00", -- $0aedd
          44766 => x"00", -- $0aede
          44767 => x"00", -- $0aedf
          44768 => x"00", -- $0aee0
          44769 => x"00", -- $0aee1
          44770 => x"00", -- $0aee2
          44771 => x"00", -- $0aee3
          44772 => x"00", -- $0aee4
          44773 => x"00", -- $0aee5
          44774 => x"00", -- $0aee6
          44775 => x"00", -- $0aee7
          44776 => x"00", -- $0aee8
          44777 => x"00", -- $0aee9
          44778 => x"00", -- $0aeea
          44779 => x"00", -- $0aeeb
          44780 => x"00", -- $0aeec
          44781 => x"00", -- $0aeed
          44782 => x"00", -- $0aeee
          44783 => x"00", -- $0aeef
          44784 => x"00", -- $0aef0
          44785 => x"00", -- $0aef1
          44786 => x"00", -- $0aef2
          44787 => x"00", -- $0aef3
          44788 => x"00", -- $0aef4
          44789 => x"00", -- $0aef5
          44790 => x"00", -- $0aef6
          44791 => x"00", -- $0aef7
          44792 => x"00", -- $0aef8
          44793 => x"00", -- $0aef9
          44794 => x"00", -- $0aefa
          44795 => x"00", -- $0aefb
          44796 => x"00", -- $0aefc
          44797 => x"00", -- $0aefd
          44798 => x"00", -- $0aefe
          44799 => x"00", -- $0aeff
          44800 => x"00", -- $0af00
          44801 => x"00", -- $0af01
          44802 => x"00", -- $0af02
          44803 => x"00", -- $0af03
          44804 => x"00", -- $0af04
          44805 => x"00", -- $0af05
          44806 => x"00", -- $0af06
          44807 => x"00", -- $0af07
          44808 => x"00", -- $0af08
          44809 => x"00", -- $0af09
          44810 => x"00", -- $0af0a
          44811 => x"00", -- $0af0b
          44812 => x"00", -- $0af0c
          44813 => x"00", -- $0af0d
          44814 => x"00", -- $0af0e
          44815 => x"00", -- $0af0f
          44816 => x"00", -- $0af10
          44817 => x"00", -- $0af11
          44818 => x"00", -- $0af12
          44819 => x"00", -- $0af13
          44820 => x"00", -- $0af14
          44821 => x"00", -- $0af15
          44822 => x"00", -- $0af16
          44823 => x"00", -- $0af17
          44824 => x"00", -- $0af18
          44825 => x"00", -- $0af19
          44826 => x"00", -- $0af1a
          44827 => x"00", -- $0af1b
          44828 => x"00", -- $0af1c
          44829 => x"00", -- $0af1d
          44830 => x"00", -- $0af1e
          44831 => x"00", -- $0af1f
          44832 => x"00", -- $0af20
          44833 => x"00", -- $0af21
          44834 => x"00", -- $0af22
          44835 => x"00", -- $0af23
          44836 => x"00", -- $0af24
          44837 => x"00", -- $0af25
          44838 => x"00", -- $0af26
          44839 => x"00", -- $0af27
          44840 => x"00", -- $0af28
          44841 => x"00", -- $0af29
          44842 => x"00", -- $0af2a
          44843 => x"00", -- $0af2b
          44844 => x"00", -- $0af2c
          44845 => x"00", -- $0af2d
          44846 => x"00", -- $0af2e
          44847 => x"00", -- $0af2f
          44848 => x"00", -- $0af30
          44849 => x"00", -- $0af31
          44850 => x"00", -- $0af32
          44851 => x"00", -- $0af33
          44852 => x"00", -- $0af34
          44853 => x"00", -- $0af35
          44854 => x"00", -- $0af36
          44855 => x"00", -- $0af37
          44856 => x"00", -- $0af38
          44857 => x"00", -- $0af39
          44858 => x"00", -- $0af3a
          44859 => x"00", -- $0af3b
          44860 => x"00", -- $0af3c
          44861 => x"00", -- $0af3d
          44862 => x"00", -- $0af3e
          44863 => x"00", -- $0af3f
          44864 => x"00", -- $0af40
          44865 => x"00", -- $0af41
          44866 => x"00", -- $0af42
          44867 => x"00", -- $0af43
          44868 => x"00", -- $0af44
          44869 => x"00", -- $0af45
          44870 => x"00", -- $0af46
          44871 => x"00", -- $0af47
          44872 => x"00", -- $0af48
          44873 => x"00", -- $0af49
          44874 => x"00", -- $0af4a
          44875 => x"00", -- $0af4b
          44876 => x"00", -- $0af4c
          44877 => x"00", -- $0af4d
          44878 => x"00", -- $0af4e
          44879 => x"00", -- $0af4f
          44880 => x"00", -- $0af50
          44881 => x"00", -- $0af51
          44882 => x"00", -- $0af52
          44883 => x"00", -- $0af53
          44884 => x"00", -- $0af54
          44885 => x"00", -- $0af55
          44886 => x"00", -- $0af56
          44887 => x"00", -- $0af57
          44888 => x"00", -- $0af58
          44889 => x"00", -- $0af59
          44890 => x"00", -- $0af5a
          44891 => x"00", -- $0af5b
          44892 => x"00", -- $0af5c
          44893 => x"00", -- $0af5d
          44894 => x"00", -- $0af5e
          44895 => x"00", -- $0af5f
          44896 => x"00", -- $0af60
          44897 => x"00", -- $0af61
          44898 => x"00", -- $0af62
          44899 => x"00", -- $0af63
          44900 => x"00", -- $0af64
          44901 => x"00", -- $0af65
          44902 => x"00", -- $0af66
          44903 => x"00", -- $0af67
          44904 => x"00", -- $0af68
          44905 => x"00", -- $0af69
          44906 => x"00", -- $0af6a
          44907 => x"00", -- $0af6b
          44908 => x"00", -- $0af6c
          44909 => x"00", -- $0af6d
          44910 => x"00", -- $0af6e
          44911 => x"00", -- $0af6f
          44912 => x"00", -- $0af70
          44913 => x"00", -- $0af71
          44914 => x"00", -- $0af72
          44915 => x"00", -- $0af73
          44916 => x"00", -- $0af74
          44917 => x"00", -- $0af75
          44918 => x"00", -- $0af76
          44919 => x"00", -- $0af77
          44920 => x"00", -- $0af78
          44921 => x"00", -- $0af79
          44922 => x"00", -- $0af7a
          44923 => x"00", -- $0af7b
          44924 => x"00", -- $0af7c
          44925 => x"00", -- $0af7d
          44926 => x"00", -- $0af7e
          44927 => x"00", -- $0af7f
          44928 => x"00", -- $0af80
          44929 => x"00", -- $0af81
          44930 => x"00", -- $0af82
          44931 => x"00", -- $0af83
          44932 => x"00", -- $0af84
          44933 => x"00", -- $0af85
          44934 => x"00", -- $0af86
          44935 => x"00", -- $0af87
          44936 => x"00", -- $0af88
          44937 => x"00", -- $0af89
          44938 => x"00", -- $0af8a
          44939 => x"00", -- $0af8b
          44940 => x"00", -- $0af8c
          44941 => x"00", -- $0af8d
          44942 => x"00", -- $0af8e
          44943 => x"00", -- $0af8f
          44944 => x"00", -- $0af90
          44945 => x"00", -- $0af91
          44946 => x"00", -- $0af92
          44947 => x"00", -- $0af93
          44948 => x"00", -- $0af94
          44949 => x"00", -- $0af95
          44950 => x"00", -- $0af96
          44951 => x"00", -- $0af97
          44952 => x"00", -- $0af98
          44953 => x"00", -- $0af99
          44954 => x"00", -- $0af9a
          44955 => x"00", -- $0af9b
          44956 => x"00", -- $0af9c
          44957 => x"00", -- $0af9d
          44958 => x"00", -- $0af9e
          44959 => x"00", -- $0af9f
          44960 => x"00", -- $0afa0
          44961 => x"00", -- $0afa1
          44962 => x"00", -- $0afa2
          44963 => x"00", -- $0afa3
          44964 => x"00", -- $0afa4
          44965 => x"00", -- $0afa5
          44966 => x"00", -- $0afa6
          44967 => x"00", -- $0afa7
          44968 => x"00", -- $0afa8
          44969 => x"00", -- $0afa9
          44970 => x"00", -- $0afaa
          44971 => x"00", -- $0afab
          44972 => x"00", -- $0afac
          44973 => x"00", -- $0afad
          44974 => x"00", -- $0afae
          44975 => x"00", -- $0afaf
          44976 => x"00", -- $0afb0
          44977 => x"00", -- $0afb1
          44978 => x"00", -- $0afb2
          44979 => x"00", -- $0afb3
          44980 => x"00", -- $0afb4
          44981 => x"00", -- $0afb5
          44982 => x"00", -- $0afb6
          44983 => x"00", -- $0afb7
          44984 => x"00", -- $0afb8
          44985 => x"00", -- $0afb9
          44986 => x"00", -- $0afba
          44987 => x"00", -- $0afbb
          44988 => x"00", -- $0afbc
          44989 => x"00", -- $0afbd
          44990 => x"00", -- $0afbe
          44991 => x"00", -- $0afbf
          44992 => x"00", -- $0afc0
          44993 => x"00", -- $0afc1
          44994 => x"00", -- $0afc2
          44995 => x"00", -- $0afc3
          44996 => x"00", -- $0afc4
          44997 => x"00", -- $0afc5
          44998 => x"00", -- $0afc6
          44999 => x"00", -- $0afc7
          45000 => x"00", -- $0afc8
          45001 => x"00", -- $0afc9
          45002 => x"00", -- $0afca
          45003 => x"00", -- $0afcb
          45004 => x"00", -- $0afcc
          45005 => x"00", -- $0afcd
          45006 => x"00", -- $0afce
          45007 => x"00", -- $0afcf
          45008 => x"00", -- $0afd0
          45009 => x"00", -- $0afd1
          45010 => x"00", -- $0afd2
          45011 => x"00", -- $0afd3
          45012 => x"00", -- $0afd4
          45013 => x"00", -- $0afd5
          45014 => x"00", -- $0afd6
          45015 => x"00", -- $0afd7
          45016 => x"00", -- $0afd8
          45017 => x"00", -- $0afd9
          45018 => x"00", -- $0afda
          45019 => x"00", -- $0afdb
          45020 => x"00", -- $0afdc
          45021 => x"00", -- $0afdd
          45022 => x"00", -- $0afde
          45023 => x"00", -- $0afdf
          45024 => x"00", -- $0afe0
          45025 => x"00", -- $0afe1
          45026 => x"00", -- $0afe2
          45027 => x"00", -- $0afe3
          45028 => x"00", -- $0afe4
          45029 => x"00", -- $0afe5
          45030 => x"00", -- $0afe6
          45031 => x"00", -- $0afe7
          45032 => x"00", -- $0afe8
          45033 => x"00", -- $0afe9
          45034 => x"00", -- $0afea
          45035 => x"00", -- $0afeb
          45036 => x"00", -- $0afec
          45037 => x"00", -- $0afed
          45038 => x"00", -- $0afee
          45039 => x"00", -- $0afef
          45040 => x"00", -- $0aff0
          45041 => x"00", -- $0aff1
          45042 => x"00", -- $0aff2
          45043 => x"00", -- $0aff3
          45044 => x"00", -- $0aff4
          45045 => x"00", -- $0aff5
          45046 => x"00", -- $0aff6
          45047 => x"00", -- $0aff7
          45048 => x"00", -- $0aff8
          45049 => x"00", -- $0aff9
          45050 => x"00", -- $0affa
          45051 => x"00", -- $0affb
          45052 => x"00", -- $0affc
          45053 => x"00", -- $0affd
          45054 => x"00", -- $0affe
          45055 => x"00", -- $0afff
          45056 => x"00", -- $0b000
          45057 => x"00", -- $0b001
          45058 => x"00", -- $0b002
          45059 => x"00", -- $0b003
          45060 => x"00", -- $0b004
          45061 => x"00", -- $0b005
          45062 => x"00", -- $0b006
          45063 => x"00", -- $0b007
          45064 => x"00", -- $0b008
          45065 => x"00", -- $0b009
          45066 => x"00", -- $0b00a
          45067 => x"00", -- $0b00b
          45068 => x"00", -- $0b00c
          45069 => x"00", -- $0b00d
          45070 => x"00", -- $0b00e
          45071 => x"00", -- $0b00f
          45072 => x"00", -- $0b010
          45073 => x"00", -- $0b011
          45074 => x"00", -- $0b012
          45075 => x"00", -- $0b013
          45076 => x"00", -- $0b014
          45077 => x"00", -- $0b015
          45078 => x"00", -- $0b016
          45079 => x"00", -- $0b017
          45080 => x"00", -- $0b018
          45081 => x"00", -- $0b019
          45082 => x"00", -- $0b01a
          45083 => x"00", -- $0b01b
          45084 => x"00", -- $0b01c
          45085 => x"00", -- $0b01d
          45086 => x"00", -- $0b01e
          45087 => x"00", -- $0b01f
          45088 => x"00", -- $0b020
          45089 => x"00", -- $0b021
          45090 => x"00", -- $0b022
          45091 => x"00", -- $0b023
          45092 => x"00", -- $0b024
          45093 => x"00", -- $0b025
          45094 => x"00", -- $0b026
          45095 => x"00", -- $0b027
          45096 => x"00", -- $0b028
          45097 => x"00", -- $0b029
          45098 => x"00", -- $0b02a
          45099 => x"00", -- $0b02b
          45100 => x"00", -- $0b02c
          45101 => x"00", -- $0b02d
          45102 => x"00", -- $0b02e
          45103 => x"00", -- $0b02f
          45104 => x"00", -- $0b030
          45105 => x"00", -- $0b031
          45106 => x"00", -- $0b032
          45107 => x"00", -- $0b033
          45108 => x"00", -- $0b034
          45109 => x"00", -- $0b035
          45110 => x"00", -- $0b036
          45111 => x"00", -- $0b037
          45112 => x"00", -- $0b038
          45113 => x"00", -- $0b039
          45114 => x"00", -- $0b03a
          45115 => x"00", -- $0b03b
          45116 => x"00", -- $0b03c
          45117 => x"00", -- $0b03d
          45118 => x"00", -- $0b03e
          45119 => x"00", -- $0b03f
          45120 => x"00", -- $0b040
          45121 => x"00", -- $0b041
          45122 => x"00", -- $0b042
          45123 => x"00", -- $0b043
          45124 => x"00", -- $0b044
          45125 => x"00", -- $0b045
          45126 => x"00", -- $0b046
          45127 => x"00", -- $0b047
          45128 => x"00", -- $0b048
          45129 => x"00", -- $0b049
          45130 => x"00", -- $0b04a
          45131 => x"00", -- $0b04b
          45132 => x"00", -- $0b04c
          45133 => x"00", -- $0b04d
          45134 => x"00", -- $0b04e
          45135 => x"00", -- $0b04f
          45136 => x"00", -- $0b050
          45137 => x"00", -- $0b051
          45138 => x"00", -- $0b052
          45139 => x"00", -- $0b053
          45140 => x"00", -- $0b054
          45141 => x"00", -- $0b055
          45142 => x"00", -- $0b056
          45143 => x"00", -- $0b057
          45144 => x"00", -- $0b058
          45145 => x"00", -- $0b059
          45146 => x"00", -- $0b05a
          45147 => x"00", -- $0b05b
          45148 => x"00", -- $0b05c
          45149 => x"00", -- $0b05d
          45150 => x"00", -- $0b05e
          45151 => x"00", -- $0b05f
          45152 => x"00", -- $0b060
          45153 => x"00", -- $0b061
          45154 => x"00", -- $0b062
          45155 => x"00", -- $0b063
          45156 => x"00", -- $0b064
          45157 => x"00", -- $0b065
          45158 => x"00", -- $0b066
          45159 => x"00", -- $0b067
          45160 => x"00", -- $0b068
          45161 => x"00", -- $0b069
          45162 => x"00", -- $0b06a
          45163 => x"00", -- $0b06b
          45164 => x"00", -- $0b06c
          45165 => x"00", -- $0b06d
          45166 => x"00", -- $0b06e
          45167 => x"00", -- $0b06f
          45168 => x"00", -- $0b070
          45169 => x"00", -- $0b071
          45170 => x"00", -- $0b072
          45171 => x"00", -- $0b073
          45172 => x"00", -- $0b074
          45173 => x"00", -- $0b075
          45174 => x"00", -- $0b076
          45175 => x"00", -- $0b077
          45176 => x"00", -- $0b078
          45177 => x"00", -- $0b079
          45178 => x"00", -- $0b07a
          45179 => x"00", -- $0b07b
          45180 => x"00", -- $0b07c
          45181 => x"00", -- $0b07d
          45182 => x"00", -- $0b07e
          45183 => x"00", -- $0b07f
          45184 => x"00", -- $0b080
          45185 => x"00", -- $0b081
          45186 => x"00", -- $0b082
          45187 => x"00", -- $0b083
          45188 => x"00", -- $0b084
          45189 => x"00", -- $0b085
          45190 => x"00", -- $0b086
          45191 => x"00", -- $0b087
          45192 => x"00", -- $0b088
          45193 => x"00", -- $0b089
          45194 => x"00", -- $0b08a
          45195 => x"00", -- $0b08b
          45196 => x"00", -- $0b08c
          45197 => x"00", -- $0b08d
          45198 => x"00", -- $0b08e
          45199 => x"00", -- $0b08f
          45200 => x"00", -- $0b090
          45201 => x"00", -- $0b091
          45202 => x"00", -- $0b092
          45203 => x"00", -- $0b093
          45204 => x"00", -- $0b094
          45205 => x"00", -- $0b095
          45206 => x"00", -- $0b096
          45207 => x"00", -- $0b097
          45208 => x"00", -- $0b098
          45209 => x"00", -- $0b099
          45210 => x"00", -- $0b09a
          45211 => x"00", -- $0b09b
          45212 => x"00", -- $0b09c
          45213 => x"00", -- $0b09d
          45214 => x"00", -- $0b09e
          45215 => x"00", -- $0b09f
          45216 => x"00", -- $0b0a0
          45217 => x"00", -- $0b0a1
          45218 => x"00", -- $0b0a2
          45219 => x"00", -- $0b0a3
          45220 => x"00", -- $0b0a4
          45221 => x"00", -- $0b0a5
          45222 => x"00", -- $0b0a6
          45223 => x"00", -- $0b0a7
          45224 => x"00", -- $0b0a8
          45225 => x"00", -- $0b0a9
          45226 => x"00", -- $0b0aa
          45227 => x"00", -- $0b0ab
          45228 => x"00", -- $0b0ac
          45229 => x"00", -- $0b0ad
          45230 => x"00", -- $0b0ae
          45231 => x"00", -- $0b0af
          45232 => x"00", -- $0b0b0
          45233 => x"00", -- $0b0b1
          45234 => x"00", -- $0b0b2
          45235 => x"00", -- $0b0b3
          45236 => x"00", -- $0b0b4
          45237 => x"00", -- $0b0b5
          45238 => x"00", -- $0b0b6
          45239 => x"00", -- $0b0b7
          45240 => x"00", -- $0b0b8
          45241 => x"00", -- $0b0b9
          45242 => x"00", -- $0b0ba
          45243 => x"00", -- $0b0bb
          45244 => x"00", -- $0b0bc
          45245 => x"00", -- $0b0bd
          45246 => x"00", -- $0b0be
          45247 => x"00", -- $0b0bf
          45248 => x"00", -- $0b0c0
          45249 => x"00", -- $0b0c1
          45250 => x"00", -- $0b0c2
          45251 => x"00", -- $0b0c3
          45252 => x"00", -- $0b0c4
          45253 => x"00", -- $0b0c5
          45254 => x"00", -- $0b0c6
          45255 => x"00", -- $0b0c7
          45256 => x"00", -- $0b0c8
          45257 => x"00", -- $0b0c9
          45258 => x"00", -- $0b0ca
          45259 => x"00", -- $0b0cb
          45260 => x"00", -- $0b0cc
          45261 => x"00", -- $0b0cd
          45262 => x"00", -- $0b0ce
          45263 => x"00", -- $0b0cf
          45264 => x"00", -- $0b0d0
          45265 => x"00", -- $0b0d1
          45266 => x"00", -- $0b0d2
          45267 => x"00", -- $0b0d3
          45268 => x"00", -- $0b0d4
          45269 => x"00", -- $0b0d5
          45270 => x"00", -- $0b0d6
          45271 => x"00", -- $0b0d7
          45272 => x"00", -- $0b0d8
          45273 => x"00", -- $0b0d9
          45274 => x"00", -- $0b0da
          45275 => x"00", -- $0b0db
          45276 => x"00", -- $0b0dc
          45277 => x"00", -- $0b0dd
          45278 => x"00", -- $0b0de
          45279 => x"00", -- $0b0df
          45280 => x"00", -- $0b0e0
          45281 => x"00", -- $0b0e1
          45282 => x"00", -- $0b0e2
          45283 => x"00", -- $0b0e3
          45284 => x"00", -- $0b0e4
          45285 => x"00", -- $0b0e5
          45286 => x"00", -- $0b0e6
          45287 => x"00", -- $0b0e7
          45288 => x"00", -- $0b0e8
          45289 => x"00", -- $0b0e9
          45290 => x"00", -- $0b0ea
          45291 => x"00", -- $0b0eb
          45292 => x"00", -- $0b0ec
          45293 => x"00", -- $0b0ed
          45294 => x"00", -- $0b0ee
          45295 => x"00", -- $0b0ef
          45296 => x"00", -- $0b0f0
          45297 => x"00", -- $0b0f1
          45298 => x"00", -- $0b0f2
          45299 => x"00", -- $0b0f3
          45300 => x"00", -- $0b0f4
          45301 => x"00", -- $0b0f5
          45302 => x"00", -- $0b0f6
          45303 => x"00", -- $0b0f7
          45304 => x"00", -- $0b0f8
          45305 => x"00", -- $0b0f9
          45306 => x"00", -- $0b0fa
          45307 => x"00", -- $0b0fb
          45308 => x"00", -- $0b0fc
          45309 => x"00", -- $0b0fd
          45310 => x"00", -- $0b0fe
          45311 => x"00", -- $0b0ff
          45312 => x"00", -- $0b100
          45313 => x"00", -- $0b101
          45314 => x"00", -- $0b102
          45315 => x"00", -- $0b103
          45316 => x"00", -- $0b104
          45317 => x"00", -- $0b105
          45318 => x"00", -- $0b106
          45319 => x"00", -- $0b107
          45320 => x"00", -- $0b108
          45321 => x"00", -- $0b109
          45322 => x"00", -- $0b10a
          45323 => x"00", -- $0b10b
          45324 => x"00", -- $0b10c
          45325 => x"00", -- $0b10d
          45326 => x"00", -- $0b10e
          45327 => x"00", -- $0b10f
          45328 => x"00", -- $0b110
          45329 => x"00", -- $0b111
          45330 => x"00", -- $0b112
          45331 => x"00", -- $0b113
          45332 => x"00", -- $0b114
          45333 => x"00", -- $0b115
          45334 => x"00", -- $0b116
          45335 => x"00", -- $0b117
          45336 => x"00", -- $0b118
          45337 => x"00", -- $0b119
          45338 => x"00", -- $0b11a
          45339 => x"00", -- $0b11b
          45340 => x"00", -- $0b11c
          45341 => x"00", -- $0b11d
          45342 => x"00", -- $0b11e
          45343 => x"00", -- $0b11f
          45344 => x"00", -- $0b120
          45345 => x"00", -- $0b121
          45346 => x"00", -- $0b122
          45347 => x"00", -- $0b123
          45348 => x"00", -- $0b124
          45349 => x"00", -- $0b125
          45350 => x"00", -- $0b126
          45351 => x"00", -- $0b127
          45352 => x"00", -- $0b128
          45353 => x"00", -- $0b129
          45354 => x"00", -- $0b12a
          45355 => x"00", -- $0b12b
          45356 => x"00", -- $0b12c
          45357 => x"00", -- $0b12d
          45358 => x"00", -- $0b12e
          45359 => x"00", -- $0b12f
          45360 => x"00", -- $0b130
          45361 => x"00", -- $0b131
          45362 => x"00", -- $0b132
          45363 => x"00", -- $0b133
          45364 => x"00", -- $0b134
          45365 => x"00", -- $0b135
          45366 => x"00", -- $0b136
          45367 => x"00", -- $0b137
          45368 => x"00", -- $0b138
          45369 => x"00", -- $0b139
          45370 => x"00", -- $0b13a
          45371 => x"00", -- $0b13b
          45372 => x"00", -- $0b13c
          45373 => x"00", -- $0b13d
          45374 => x"00", -- $0b13e
          45375 => x"00", -- $0b13f
          45376 => x"00", -- $0b140
          45377 => x"00", -- $0b141
          45378 => x"00", -- $0b142
          45379 => x"00", -- $0b143
          45380 => x"00", -- $0b144
          45381 => x"00", -- $0b145
          45382 => x"00", -- $0b146
          45383 => x"00", -- $0b147
          45384 => x"00", -- $0b148
          45385 => x"00", -- $0b149
          45386 => x"00", -- $0b14a
          45387 => x"00", -- $0b14b
          45388 => x"00", -- $0b14c
          45389 => x"00", -- $0b14d
          45390 => x"00", -- $0b14e
          45391 => x"00", -- $0b14f
          45392 => x"00", -- $0b150
          45393 => x"00", -- $0b151
          45394 => x"00", -- $0b152
          45395 => x"00", -- $0b153
          45396 => x"00", -- $0b154
          45397 => x"00", -- $0b155
          45398 => x"00", -- $0b156
          45399 => x"00", -- $0b157
          45400 => x"00", -- $0b158
          45401 => x"00", -- $0b159
          45402 => x"00", -- $0b15a
          45403 => x"00", -- $0b15b
          45404 => x"00", -- $0b15c
          45405 => x"00", -- $0b15d
          45406 => x"00", -- $0b15e
          45407 => x"00", -- $0b15f
          45408 => x"00", -- $0b160
          45409 => x"00", -- $0b161
          45410 => x"00", -- $0b162
          45411 => x"00", -- $0b163
          45412 => x"00", -- $0b164
          45413 => x"00", -- $0b165
          45414 => x"00", -- $0b166
          45415 => x"00", -- $0b167
          45416 => x"00", -- $0b168
          45417 => x"00", -- $0b169
          45418 => x"00", -- $0b16a
          45419 => x"00", -- $0b16b
          45420 => x"00", -- $0b16c
          45421 => x"00", -- $0b16d
          45422 => x"00", -- $0b16e
          45423 => x"00", -- $0b16f
          45424 => x"00", -- $0b170
          45425 => x"00", -- $0b171
          45426 => x"00", -- $0b172
          45427 => x"00", -- $0b173
          45428 => x"00", -- $0b174
          45429 => x"00", -- $0b175
          45430 => x"00", -- $0b176
          45431 => x"00", -- $0b177
          45432 => x"00", -- $0b178
          45433 => x"00", -- $0b179
          45434 => x"00", -- $0b17a
          45435 => x"00", -- $0b17b
          45436 => x"00", -- $0b17c
          45437 => x"00", -- $0b17d
          45438 => x"00", -- $0b17e
          45439 => x"00", -- $0b17f
          45440 => x"00", -- $0b180
          45441 => x"00", -- $0b181
          45442 => x"00", -- $0b182
          45443 => x"00", -- $0b183
          45444 => x"00", -- $0b184
          45445 => x"00", -- $0b185
          45446 => x"00", -- $0b186
          45447 => x"00", -- $0b187
          45448 => x"00", -- $0b188
          45449 => x"00", -- $0b189
          45450 => x"00", -- $0b18a
          45451 => x"00", -- $0b18b
          45452 => x"00", -- $0b18c
          45453 => x"00", -- $0b18d
          45454 => x"00", -- $0b18e
          45455 => x"00", -- $0b18f
          45456 => x"00", -- $0b190
          45457 => x"00", -- $0b191
          45458 => x"00", -- $0b192
          45459 => x"00", -- $0b193
          45460 => x"00", -- $0b194
          45461 => x"00", -- $0b195
          45462 => x"00", -- $0b196
          45463 => x"00", -- $0b197
          45464 => x"00", -- $0b198
          45465 => x"00", -- $0b199
          45466 => x"00", -- $0b19a
          45467 => x"00", -- $0b19b
          45468 => x"00", -- $0b19c
          45469 => x"00", -- $0b19d
          45470 => x"00", -- $0b19e
          45471 => x"00", -- $0b19f
          45472 => x"00", -- $0b1a0
          45473 => x"00", -- $0b1a1
          45474 => x"00", -- $0b1a2
          45475 => x"00", -- $0b1a3
          45476 => x"00", -- $0b1a4
          45477 => x"00", -- $0b1a5
          45478 => x"00", -- $0b1a6
          45479 => x"00", -- $0b1a7
          45480 => x"00", -- $0b1a8
          45481 => x"00", -- $0b1a9
          45482 => x"00", -- $0b1aa
          45483 => x"00", -- $0b1ab
          45484 => x"00", -- $0b1ac
          45485 => x"00", -- $0b1ad
          45486 => x"00", -- $0b1ae
          45487 => x"00", -- $0b1af
          45488 => x"00", -- $0b1b0
          45489 => x"00", -- $0b1b1
          45490 => x"00", -- $0b1b2
          45491 => x"00", -- $0b1b3
          45492 => x"00", -- $0b1b4
          45493 => x"00", -- $0b1b5
          45494 => x"00", -- $0b1b6
          45495 => x"00", -- $0b1b7
          45496 => x"00", -- $0b1b8
          45497 => x"00", -- $0b1b9
          45498 => x"00", -- $0b1ba
          45499 => x"00", -- $0b1bb
          45500 => x"00", -- $0b1bc
          45501 => x"00", -- $0b1bd
          45502 => x"00", -- $0b1be
          45503 => x"00", -- $0b1bf
          45504 => x"00", -- $0b1c0
          45505 => x"00", -- $0b1c1
          45506 => x"00", -- $0b1c2
          45507 => x"00", -- $0b1c3
          45508 => x"00", -- $0b1c4
          45509 => x"00", -- $0b1c5
          45510 => x"00", -- $0b1c6
          45511 => x"00", -- $0b1c7
          45512 => x"00", -- $0b1c8
          45513 => x"00", -- $0b1c9
          45514 => x"00", -- $0b1ca
          45515 => x"00", -- $0b1cb
          45516 => x"00", -- $0b1cc
          45517 => x"00", -- $0b1cd
          45518 => x"00", -- $0b1ce
          45519 => x"00", -- $0b1cf
          45520 => x"00", -- $0b1d0
          45521 => x"00", -- $0b1d1
          45522 => x"00", -- $0b1d2
          45523 => x"00", -- $0b1d3
          45524 => x"00", -- $0b1d4
          45525 => x"00", -- $0b1d5
          45526 => x"00", -- $0b1d6
          45527 => x"00", -- $0b1d7
          45528 => x"00", -- $0b1d8
          45529 => x"00", -- $0b1d9
          45530 => x"00", -- $0b1da
          45531 => x"00", -- $0b1db
          45532 => x"00", -- $0b1dc
          45533 => x"00", -- $0b1dd
          45534 => x"00", -- $0b1de
          45535 => x"00", -- $0b1df
          45536 => x"00", -- $0b1e0
          45537 => x"00", -- $0b1e1
          45538 => x"00", -- $0b1e2
          45539 => x"00", -- $0b1e3
          45540 => x"00", -- $0b1e4
          45541 => x"00", -- $0b1e5
          45542 => x"00", -- $0b1e6
          45543 => x"00", -- $0b1e7
          45544 => x"00", -- $0b1e8
          45545 => x"00", -- $0b1e9
          45546 => x"00", -- $0b1ea
          45547 => x"00", -- $0b1eb
          45548 => x"00", -- $0b1ec
          45549 => x"00", -- $0b1ed
          45550 => x"00", -- $0b1ee
          45551 => x"00", -- $0b1ef
          45552 => x"00", -- $0b1f0
          45553 => x"00", -- $0b1f1
          45554 => x"00", -- $0b1f2
          45555 => x"00", -- $0b1f3
          45556 => x"00", -- $0b1f4
          45557 => x"00", -- $0b1f5
          45558 => x"00", -- $0b1f6
          45559 => x"00", -- $0b1f7
          45560 => x"00", -- $0b1f8
          45561 => x"00", -- $0b1f9
          45562 => x"00", -- $0b1fa
          45563 => x"00", -- $0b1fb
          45564 => x"00", -- $0b1fc
          45565 => x"00", -- $0b1fd
          45566 => x"00", -- $0b1fe
          45567 => x"00", -- $0b1ff
          45568 => x"00", -- $0b200
          45569 => x"00", -- $0b201
          45570 => x"00", -- $0b202
          45571 => x"00", -- $0b203
          45572 => x"00", -- $0b204
          45573 => x"00", -- $0b205
          45574 => x"00", -- $0b206
          45575 => x"00", -- $0b207
          45576 => x"00", -- $0b208
          45577 => x"00", -- $0b209
          45578 => x"00", -- $0b20a
          45579 => x"00", -- $0b20b
          45580 => x"00", -- $0b20c
          45581 => x"00", -- $0b20d
          45582 => x"00", -- $0b20e
          45583 => x"00", -- $0b20f
          45584 => x"00", -- $0b210
          45585 => x"00", -- $0b211
          45586 => x"00", -- $0b212
          45587 => x"00", -- $0b213
          45588 => x"00", -- $0b214
          45589 => x"00", -- $0b215
          45590 => x"00", -- $0b216
          45591 => x"00", -- $0b217
          45592 => x"00", -- $0b218
          45593 => x"00", -- $0b219
          45594 => x"00", -- $0b21a
          45595 => x"00", -- $0b21b
          45596 => x"00", -- $0b21c
          45597 => x"00", -- $0b21d
          45598 => x"00", -- $0b21e
          45599 => x"00", -- $0b21f
          45600 => x"00", -- $0b220
          45601 => x"00", -- $0b221
          45602 => x"00", -- $0b222
          45603 => x"00", -- $0b223
          45604 => x"00", -- $0b224
          45605 => x"00", -- $0b225
          45606 => x"00", -- $0b226
          45607 => x"00", -- $0b227
          45608 => x"00", -- $0b228
          45609 => x"00", -- $0b229
          45610 => x"00", -- $0b22a
          45611 => x"00", -- $0b22b
          45612 => x"00", -- $0b22c
          45613 => x"00", -- $0b22d
          45614 => x"00", -- $0b22e
          45615 => x"00", -- $0b22f
          45616 => x"00", -- $0b230
          45617 => x"00", -- $0b231
          45618 => x"00", -- $0b232
          45619 => x"00", -- $0b233
          45620 => x"00", -- $0b234
          45621 => x"00", -- $0b235
          45622 => x"00", -- $0b236
          45623 => x"00", -- $0b237
          45624 => x"00", -- $0b238
          45625 => x"00", -- $0b239
          45626 => x"00", -- $0b23a
          45627 => x"00", -- $0b23b
          45628 => x"00", -- $0b23c
          45629 => x"00", -- $0b23d
          45630 => x"00", -- $0b23e
          45631 => x"00", -- $0b23f
          45632 => x"00", -- $0b240
          45633 => x"00", -- $0b241
          45634 => x"00", -- $0b242
          45635 => x"00", -- $0b243
          45636 => x"00", -- $0b244
          45637 => x"00", -- $0b245
          45638 => x"00", -- $0b246
          45639 => x"00", -- $0b247
          45640 => x"00", -- $0b248
          45641 => x"00", -- $0b249
          45642 => x"00", -- $0b24a
          45643 => x"00", -- $0b24b
          45644 => x"00", -- $0b24c
          45645 => x"00", -- $0b24d
          45646 => x"00", -- $0b24e
          45647 => x"00", -- $0b24f
          45648 => x"00", -- $0b250
          45649 => x"00", -- $0b251
          45650 => x"00", -- $0b252
          45651 => x"00", -- $0b253
          45652 => x"00", -- $0b254
          45653 => x"00", -- $0b255
          45654 => x"00", -- $0b256
          45655 => x"00", -- $0b257
          45656 => x"00", -- $0b258
          45657 => x"00", -- $0b259
          45658 => x"00", -- $0b25a
          45659 => x"00", -- $0b25b
          45660 => x"00", -- $0b25c
          45661 => x"00", -- $0b25d
          45662 => x"00", -- $0b25e
          45663 => x"00", -- $0b25f
          45664 => x"00", -- $0b260
          45665 => x"00", -- $0b261
          45666 => x"00", -- $0b262
          45667 => x"00", -- $0b263
          45668 => x"00", -- $0b264
          45669 => x"00", -- $0b265
          45670 => x"00", -- $0b266
          45671 => x"00", -- $0b267
          45672 => x"00", -- $0b268
          45673 => x"00", -- $0b269
          45674 => x"00", -- $0b26a
          45675 => x"00", -- $0b26b
          45676 => x"00", -- $0b26c
          45677 => x"00", -- $0b26d
          45678 => x"00", -- $0b26e
          45679 => x"00", -- $0b26f
          45680 => x"00", -- $0b270
          45681 => x"00", -- $0b271
          45682 => x"00", -- $0b272
          45683 => x"00", -- $0b273
          45684 => x"00", -- $0b274
          45685 => x"00", -- $0b275
          45686 => x"00", -- $0b276
          45687 => x"00", -- $0b277
          45688 => x"00", -- $0b278
          45689 => x"00", -- $0b279
          45690 => x"00", -- $0b27a
          45691 => x"00", -- $0b27b
          45692 => x"00", -- $0b27c
          45693 => x"00", -- $0b27d
          45694 => x"00", -- $0b27e
          45695 => x"00", -- $0b27f
          45696 => x"00", -- $0b280
          45697 => x"00", -- $0b281
          45698 => x"00", -- $0b282
          45699 => x"00", -- $0b283
          45700 => x"00", -- $0b284
          45701 => x"00", -- $0b285
          45702 => x"00", -- $0b286
          45703 => x"00", -- $0b287
          45704 => x"00", -- $0b288
          45705 => x"00", -- $0b289
          45706 => x"00", -- $0b28a
          45707 => x"00", -- $0b28b
          45708 => x"00", -- $0b28c
          45709 => x"00", -- $0b28d
          45710 => x"00", -- $0b28e
          45711 => x"00", -- $0b28f
          45712 => x"00", -- $0b290
          45713 => x"00", -- $0b291
          45714 => x"00", -- $0b292
          45715 => x"00", -- $0b293
          45716 => x"00", -- $0b294
          45717 => x"00", -- $0b295
          45718 => x"00", -- $0b296
          45719 => x"00", -- $0b297
          45720 => x"00", -- $0b298
          45721 => x"00", -- $0b299
          45722 => x"00", -- $0b29a
          45723 => x"00", -- $0b29b
          45724 => x"00", -- $0b29c
          45725 => x"00", -- $0b29d
          45726 => x"00", -- $0b29e
          45727 => x"00", -- $0b29f
          45728 => x"00", -- $0b2a0
          45729 => x"00", -- $0b2a1
          45730 => x"00", -- $0b2a2
          45731 => x"00", -- $0b2a3
          45732 => x"00", -- $0b2a4
          45733 => x"00", -- $0b2a5
          45734 => x"00", -- $0b2a6
          45735 => x"00", -- $0b2a7
          45736 => x"00", -- $0b2a8
          45737 => x"00", -- $0b2a9
          45738 => x"00", -- $0b2aa
          45739 => x"00", -- $0b2ab
          45740 => x"00", -- $0b2ac
          45741 => x"00", -- $0b2ad
          45742 => x"00", -- $0b2ae
          45743 => x"00", -- $0b2af
          45744 => x"00", -- $0b2b0
          45745 => x"00", -- $0b2b1
          45746 => x"00", -- $0b2b2
          45747 => x"00", -- $0b2b3
          45748 => x"00", -- $0b2b4
          45749 => x"00", -- $0b2b5
          45750 => x"00", -- $0b2b6
          45751 => x"00", -- $0b2b7
          45752 => x"00", -- $0b2b8
          45753 => x"00", -- $0b2b9
          45754 => x"00", -- $0b2ba
          45755 => x"00", -- $0b2bb
          45756 => x"00", -- $0b2bc
          45757 => x"00", -- $0b2bd
          45758 => x"00", -- $0b2be
          45759 => x"00", -- $0b2bf
          45760 => x"00", -- $0b2c0
          45761 => x"00", -- $0b2c1
          45762 => x"00", -- $0b2c2
          45763 => x"00", -- $0b2c3
          45764 => x"00", -- $0b2c4
          45765 => x"00", -- $0b2c5
          45766 => x"00", -- $0b2c6
          45767 => x"00", -- $0b2c7
          45768 => x"00", -- $0b2c8
          45769 => x"00", -- $0b2c9
          45770 => x"00", -- $0b2ca
          45771 => x"00", -- $0b2cb
          45772 => x"00", -- $0b2cc
          45773 => x"00", -- $0b2cd
          45774 => x"00", -- $0b2ce
          45775 => x"00", -- $0b2cf
          45776 => x"00", -- $0b2d0
          45777 => x"00", -- $0b2d1
          45778 => x"00", -- $0b2d2
          45779 => x"00", -- $0b2d3
          45780 => x"00", -- $0b2d4
          45781 => x"00", -- $0b2d5
          45782 => x"00", -- $0b2d6
          45783 => x"00", -- $0b2d7
          45784 => x"00", -- $0b2d8
          45785 => x"00", -- $0b2d9
          45786 => x"00", -- $0b2da
          45787 => x"00", -- $0b2db
          45788 => x"00", -- $0b2dc
          45789 => x"00", -- $0b2dd
          45790 => x"00", -- $0b2de
          45791 => x"00", -- $0b2df
          45792 => x"00", -- $0b2e0
          45793 => x"00", -- $0b2e1
          45794 => x"00", -- $0b2e2
          45795 => x"00", -- $0b2e3
          45796 => x"00", -- $0b2e4
          45797 => x"00", -- $0b2e5
          45798 => x"00", -- $0b2e6
          45799 => x"00", -- $0b2e7
          45800 => x"00", -- $0b2e8
          45801 => x"00", -- $0b2e9
          45802 => x"00", -- $0b2ea
          45803 => x"00", -- $0b2eb
          45804 => x"00", -- $0b2ec
          45805 => x"00", -- $0b2ed
          45806 => x"00", -- $0b2ee
          45807 => x"00", -- $0b2ef
          45808 => x"00", -- $0b2f0
          45809 => x"00", -- $0b2f1
          45810 => x"00", -- $0b2f2
          45811 => x"00", -- $0b2f3
          45812 => x"00", -- $0b2f4
          45813 => x"00", -- $0b2f5
          45814 => x"00", -- $0b2f6
          45815 => x"00", -- $0b2f7
          45816 => x"00", -- $0b2f8
          45817 => x"00", -- $0b2f9
          45818 => x"00", -- $0b2fa
          45819 => x"00", -- $0b2fb
          45820 => x"00", -- $0b2fc
          45821 => x"00", -- $0b2fd
          45822 => x"00", -- $0b2fe
          45823 => x"00", -- $0b2ff
          45824 => x"00", -- $0b300
          45825 => x"00", -- $0b301
          45826 => x"00", -- $0b302
          45827 => x"00", -- $0b303
          45828 => x"00", -- $0b304
          45829 => x"00", -- $0b305
          45830 => x"00", -- $0b306
          45831 => x"00", -- $0b307
          45832 => x"00", -- $0b308
          45833 => x"00", -- $0b309
          45834 => x"00", -- $0b30a
          45835 => x"00", -- $0b30b
          45836 => x"00", -- $0b30c
          45837 => x"00", -- $0b30d
          45838 => x"00", -- $0b30e
          45839 => x"00", -- $0b30f
          45840 => x"00", -- $0b310
          45841 => x"00", -- $0b311
          45842 => x"00", -- $0b312
          45843 => x"00", -- $0b313
          45844 => x"00", -- $0b314
          45845 => x"00", -- $0b315
          45846 => x"00", -- $0b316
          45847 => x"00", -- $0b317
          45848 => x"00", -- $0b318
          45849 => x"00", -- $0b319
          45850 => x"00", -- $0b31a
          45851 => x"00", -- $0b31b
          45852 => x"00", -- $0b31c
          45853 => x"00", -- $0b31d
          45854 => x"00", -- $0b31e
          45855 => x"00", -- $0b31f
          45856 => x"00", -- $0b320
          45857 => x"00", -- $0b321
          45858 => x"00", -- $0b322
          45859 => x"00", -- $0b323
          45860 => x"00", -- $0b324
          45861 => x"00", -- $0b325
          45862 => x"00", -- $0b326
          45863 => x"00", -- $0b327
          45864 => x"00", -- $0b328
          45865 => x"00", -- $0b329
          45866 => x"00", -- $0b32a
          45867 => x"00", -- $0b32b
          45868 => x"00", -- $0b32c
          45869 => x"00", -- $0b32d
          45870 => x"00", -- $0b32e
          45871 => x"00", -- $0b32f
          45872 => x"00", -- $0b330
          45873 => x"00", -- $0b331
          45874 => x"00", -- $0b332
          45875 => x"00", -- $0b333
          45876 => x"00", -- $0b334
          45877 => x"00", -- $0b335
          45878 => x"00", -- $0b336
          45879 => x"00", -- $0b337
          45880 => x"00", -- $0b338
          45881 => x"00", -- $0b339
          45882 => x"00", -- $0b33a
          45883 => x"00", -- $0b33b
          45884 => x"00", -- $0b33c
          45885 => x"00", -- $0b33d
          45886 => x"00", -- $0b33e
          45887 => x"00", -- $0b33f
          45888 => x"00", -- $0b340
          45889 => x"00", -- $0b341
          45890 => x"00", -- $0b342
          45891 => x"00", -- $0b343
          45892 => x"00", -- $0b344
          45893 => x"00", -- $0b345
          45894 => x"00", -- $0b346
          45895 => x"00", -- $0b347
          45896 => x"00", -- $0b348
          45897 => x"00", -- $0b349
          45898 => x"00", -- $0b34a
          45899 => x"00", -- $0b34b
          45900 => x"00", -- $0b34c
          45901 => x"00", -- $0b34d
          45902 => x"00", -- $0b34e
          45903 => x"00", -- $0b34f
          45904 => x"00", -- $0b350
          45905 => x"00", -- $0b351
          45906 => x"00", -- $0b352
          45907 => x"00", -- $0b353
          45908 => x"00", -- $0b354
          45909 => x"00", -- $0b355
          45910 => x"00", -- $0b356
          45911 => x"00", -- $0b357
          45912 => x"00", -- $0b358
          45913 => x"00", -- $0b359
          45914 => x"00", -- $0b35a
          45915 => x"00", -- $0b35b
          45916 => x"00", -- $0b35c
          45917 => x"00", -- $0b35d
          45918 => x"00", -- $0b35e
          45919 => x"00", -- $0b35f
          45920 => x"00", -- $0b360
          45921 => x"00", -- $0b361
          45922 => x"00", -- $0b362
          45923 => x"00", -- $0b363
          45924 => x"00", -- $0b364
          45925 => x"00", -- $0b365
          45926 => x"00", -- $0b366
          45927 => x"00", -- $0b367
          45928 => x"00", -- $0b368
          45929 => x"00", -- $0b369
          45930 => x"00", -- $0b36a
          45931 => x"00", -- $0b36b
          45932 => x"00", -- $0b36c
          45933 => x"00", -- $0b36d
          45934 => x"00", -- $0b36e
          45935 => x"00", -- $0b36f
          45936 => x"00", -- $0b370
          45937 => x"00", -- $0b371
          45938 => x"00", -- $0b372
          45939 => x"00", -- $0b373
          45940 => x"00", -- $0b374
          45941 => x"00", -- $0b375
          45942 => x"00", -- $0b376
          45943 => x"00", -- $0b377
          45944 => x"00", -- $0b378
          45945 => x"00", -- $0b379
          45946 => x"00", -- $0b37a
          45947 => x"00", -- $0b37b
          45948 => x"00", -- $0b37c
          45949 => x"00", -- $0b37d
          45950 => x"00", -- $0b37e
          45951 => x"00", -- $0b37f
          45952 => x"00", -- $0b380
          45953 => x"00", -- $0b381
          45954 => x"00", -- $0b382
          45955 => x"00", -- $0b383
          45956 => x"00", -- $0b384
          45957 => x"00", -- $0b385
          45958 => x"00", -- $0b386
          45959 => x"00", -- $0b387
          45960 => x"00", -- $0b388
          45961 => x"00", -- $0b389
          45962 => x"00", -- $0b38a
          45963 => x"00", -- $0b38b
          45964 => x"00", -- $0b38c
          45965 => x"00", -- $0b38d
          45966 => x"00", -- $0b38e
          45967 => x"00", -- $0b38f
          45968 => x"00", -- $0b390
          45969 => x"00", -- $0b391
          45970 => x"00", -- $0b392
          45971 => x"00", -- $0b393
          45972 => x"00", -- $0b394
          45973 => x"00", -- $0b395
          45974 => x"00", -- $0b396
          45975 => x"00", -- $0b397
          45976 => x"00", -- $0b398
          45977 => x"00", -- $0b399
          45978 => x"00", -- $0b39a
          45979 => x"00", -- $0b39b
          45980 => x"00", -- $0b39c
          45981 => x"00", -- $0b39d
          45982 => x"00", -- $0b39e
          45983 => x"00", -- $0b39f
          45984 => x"00", -- $0b3a0
          45985 => x"00", -- $0b3a1
          45986 => x"00", -- $0b3a2
          45987 => x"00", -- $0b3a3
          45988 => x"00", -- $0b3a4
          45989 => x"00", -- $0b3a5
          45990 => x"00", -- $0b3a6
          45991 => x"00", -- $0b3a7
          45992 => x"00", -- $0b3a8
          45993 => x"00", -- $0b3a9
          45994 => x"00", -- $0b3aa
          45995 => x"00", -- $0b3ab
          45996 => x"00", -- $0b3ac
          45997 => x"00", -- $0b3ad
          45998 => x"00", -- $0b3ae
          45999 => x"00", -- $0b3af
          46000 => x"00", -- $0b3b0
          46001 => x"00", -- $0b3b1
          46002 => x"00", -- $0b3b2
          46003 => x"00", -- $0b3b3
          46004 => x"00", -- $0b3b4
          46005 => x"00", -- $0b3b5
          46006 => x"00", -- $0b3b6
          46007 => x"00", -- $0b3b7
          46008 => x"00", -- $0b3b8
          46009 => x"00", -- $0b3b9
          46010 => x"00", -- $0b3ba
          46011 => x"00", -- $0b3bb
          46012 => x"00", -- $0b3bc
          46013 => x"00", -- $0b3bd
          46014 => x"00", -- $0b3be
          46015 => x"00", -- $0b3bf
          46016 => x"00", -- $0b3c0
          46017 => x"00", -- $0b3c1
          46018 => x"00", -- $0b3c2
          46019 => x"00", -- $0b3c3
          46020 => x"00", -- $0b3c4
          46021 => x"00", -- $0b3c5
          46022 => x"00", -- $0b3c6
          46023 => x"00", -- $0b3c7
          46024 => x"00", -- $0b3c8
          46025 => x"00", -- $0b3c9
          46026 => x"00", -- $0b3ca
          46027 => x"00", -- $0b3cb
          46028 => x"00", -- $0b3cc
          46029 => x"00", -- $0b3cd
          46030 => x"00", -- $0b3ce
          46031 => x"00", -- $0b3cf
          46032 => x"00", -- $0b3d0
          46033 => x"00", -- $0b3d1
          46034 => x"00", -- $0b3d2
          46035 => x"00", -- $0b3d3
          46036 => x"00", -- $0b3d4
          46037 => x"00", -- $0b3d5
          46038 => x"00", -- $0b3d6
          46039 => x"00", -- $0b3d7
          46040 => x"00", -- $0b3d8
          46041 => x"00", -- $0b3d9
          46042 => x"00", -- $0b3da
          46043 => x"00", -- $0b3db
          46044 => x"00", -- $0b3dc
          46045 => x"00", -- $0b3dd
          46046 => x"00", -- $0b3de
          46047 => x"00", -- $0b3df
          46048 => x"00", -- $0b3e0
          46049 => x"00", -- $0b3e1
          46050 => x"00", -- $0b3e2
          46051 => x"00", -- $0b3e3
          46052 => x"00", -- $0b3e4
          46053 => x"00", -- $0b3e5
          46054 => x"00", -- $0b3e6
          46055 => x"00", -- $0b3e7
          46056 => x"00", -- $0b3e8
          46057 => x"00", -- $0b3e9
          46058 => x"00", -- $0b3ea
          46059 => x"00", -- $0b3eb
          46060 => x"00", -- $0b3ec
          46061 => x"00", -- $0b3ed
          46062 => x"00", -- $0b3ee
          46063 => x"00", -- $0b3ef
          46064 => x"00", -- $0b3f0
          46065 => x"00", -- $0b3f1
          46066 => x"00", -- $0b3f2
          46067 => x"00", -- $0b3f3
          46068 => x"00", -- $0b3f4
          46069 => x"00", -- $0b3f5
          46070 => x"00", -- $0b3f6
          46071 => x"00", -- $0b3f7
          46072 => x"00", -- $0b3f8
          46073 => x"00", -- $0b3f9
          46074 => x"00", -- $0b3fa
          46075 => x"00", -- $0b3fb
          46076 => x"00", -- $0b3fc
          46077 => x"00", -- $0b3fd
          46078 => x"00", -- $0b3fe
          46079 => x"00", -- $0b3ff
          46080 => x"00", -- $0b400
          46081 => x"00", -- $0b401
          46082 => x"00", -- $0b402
          46083 => x"00", -- $0b403
          46084 => x"00", -- $0b404
          46085 => x"00", -- $0b405
          46086 => x"00", -- $0b406
          46087 => x"00", -- $0b407
          46088 => x"00", -- $0b408
          46089 => x"00", -- $0b409
          46090 => x"00", -- $0b40a
          46091 => x"00", -- $0b40b
          46092 => x"00", -- $0b40c
          46093 => x"00", -- $0b40d
          46094 => x"00", -- $0b40e
          46095 => x"00", -- $0b40f
          46096 => x"00", -- $0b410
          46097 => x"00", -- $0b411
          46098 => x"00", -- $0b412
          46099 => x"00", -- $0b413
          46100 => x"00", -- $0b414
          46101 => x"00", -- $0b415
          46102 => x"00", -- $0b416
          46103 => x"00", -- $0b417
          46104 => x"00", -- $0b418
          46105 => x"00", -- $0b419
          46106 => x"00", -- $0b41a
          46107 => x"00", -- $0b41b
          46108 => x"00", -- $0b41c
          46109 => x"00", -- $0b41d
          46110 => x"00", -- $0b41e
          46111 => x"00", -- $0b41f
          46112 => x"00", -- $0b420
          46113 => x"00", -- $0b421
          46114 => x"00", -- $0b422
          46115 => x"00", -- $0b423
          46116 => x"00", -- $0b424
          46117 => x"00", -- $0b425
          46118 => x"00", -- $0b426
          46119 => x"00", -- $0b427
          46120 => x"00", -- $0b428
          46121 => x"00", -- $0b429
          46122 => x"00", -- $0b42a
          46123 => x"00", -- $0b42b
          46124 => x"00", -- $0b42c
          46125 => x"00", -- $0b42d
          46126 => x"00", -- $0b42e
          46127 => x"00", -- $0b42f
          46128 => x"00", -- $0b430
          46129 => x"00", -- $0b431
          46130 => x"00", -- $0b432
          46131 => x"00", -- $0b433
          46132 => x"00", -- $0b434
          46133 => x"00", -- $0b435
          46134 => x"00", -- $0b436
          46135 => x"00", -- $0b437
          46136 => x"00", -- $0b438
          46137 => x"00", -- $0b439
          46138 => x"00", -- $0b43a
          46139 => x"00", -- $0b43b
          46140 => x"00", -- $0b43c
          46141 => x"00", -- $0b43d
          46142 => x"00", -- $0b43e
          46143 => x"00", -- $0b43f
          46144 => x"00", -- $0b440
          46145 => x"00", -- $0b441
          46146 => x"00", -- $0b442
          46147 => x"00", -- $0b443
          46148 => x"00", -- $0b444
          46149 => x"00", -- $0b445
          46150 => x"00", -- $0b446
          46151 => x"00", -- $0b447
          46152 => x"00", -- $0b448
          46153 => x"00", -- $0b449
          46154 => x"00", -- $0b44a
          46155 => x"00", -- $0b44b
          46156 => x"00", -- $0b44c
          46157 => x"00", -- $0b44d
          46158 => x"00", -- $0b44e
          46159 => x"00", -- $0b44f
          46160 => x"00", -- $0b450
          46161 => x"00", -- $0b451
          46162 => x"00", -- $0b452
          46163 => x"00", -- $0b453
          46164 => x"00", -- $0b454
          46165 => x"00", -- $0b455
          46166 => x"00", -- $0b456
          46167 => x"00", -- $0b457
          46168 => x"00", -- $0b458
          46169 => x"00", -- $0b459
          46170 => x"00", -- $0b45a
          46171 => x"00", -- $0b45b
          46172 => x"00", -- $0b45c
          46173 => x"00", -- $0b45d
          46174 => x"00", -- $0b45e
          46175 => x"00", -- $0b45f
          46176 => x"00", -- $0b460
          46177 => x"00", -- $0b461
          46178 => x"00", -- $0b462
          46179 => x"00", -- $0b463
          46180 => x"00", -- $0b464
          46181 => x"00", -- $0b465
          46182 => x"00", -- $0b466
          46183 => x"00", -- $0b467
          46184 => x"00", -- $0b468
          46185 => x"00", -- $0b469
          46186 => x"00", -- $0b46a
          46187 => x"00", -- $0b46b
          46188 => x"00", -- $0b46c
          46189 => x"00", -- $0b46d
          46190 => x"00", -- $0b46e
          46191 => x"00", -- $0b46f
          46192 => x"00", -- $0b470
          46193 => x"00", -- $0b471
          46194 => x"00", -- $0b472
          46195 => x"00", -- $0b473
          46196 => x"00", -- $0b474
          46197 => x"00", -- $0b475
          46198 => x"00", -- $0b476
          46199 => x"00", -- $0b477
          46200 => x"00", -- $0b478
          46201 => x"00", -- $0b479
          46202 => x"00", -- $0b47a
          46203 => x"00", -- $0b47b
          46204 => x"00", -- $0b47c
          46205 => x"00", -- $0b47d
          46206 => x"00", -- $0b47e
          46207 => x"00", -- $0b47f
          46208 => x"00", -- $0b480
          46209 => x"00", -- $0b481
          46210 => x"00", -- $0b482
          46211 => x"00", -- $0b483
          46212 => x"00", -- $0b484
          46213 => x"00", -- $0b485
          46214 => x"00", -- $0b486
          46215 => x"00", -- $0b487
          46216 => x"00", -- $0b488
          46217 => x"00", -- $0b489
          46218 => x"00", -- $0b48a
          46219 => x"00", -- $0b48b
          46220 => x"00", -- $0b48c
          46221 => x"00", -- $0b48d
          46222 => x"00", -- $0b48e
          46223 => x"00", -- $0b48f
          46224 => x"00", -- $0b490
          46225 => x"00", -- $0b491
          46226 => x"00", -- $0b492
          46227 => x"00", -- $0b493
          46228 => x"00", -- $0b494
          46229 => x"00", -- $0b495
          46230 => x"00", -- $0b496
          46231 => x"00", -- $0b497
          46232 => x"00", -- $0b498
          46233 => x"00", -- $0b499
          46234 => x"00", -- $0b49a
          46235 => x"00", -- $0b49b
          46236 => x"00", -- $0b49c
          46237 => x"00", -- $0b49d
          46238 => x"00", -- $0b49e
          46239 => x"00", -- $0b49f
          46240 => x"00", -- $0b4a0
          46241 => x"00", -- $0b4a1
          46242 => x"00", -- $0b4a2
          46243 => x"00", -- $0b4a3
          46244 => x"00", -- $0b4a4
          46245 => x"00", -- $0b4a5
          46246 => x"00", -- $0b4a6
          46247 => x"00", -- $0b4a7
          46248 => x"00", -- $0b4a8
          46249 => x"00", -- $0b4a9
          46250 => x"00", -- $0b4aa
          46251 => x"00", -- $0b4ab
          46252 => x"00", -- $0b4ac
          46253 => x"00", -- $0b4ad
          46254 => x"00", -- $0b4ae
          46255 => x"00", -- $0b4af
          46256 => x"00", -- $0b4b0
          46257 => x"00", -- $0b4b1
          46258 => x"00", -- $0b4b2
          46259 => x"00", -- $0b4b3
          46260 => x"00", -- $0b4b4
          46261 => x"00", -- $0b4b5
          46262 => x"00", -- $0b4b6
          46263 => x"00", -- $0b4b7
          46264 => x"00", -- $0b4b8
          46265 => x"00", -- $0b4b9
          46266 => x"00", -- $0b4ba
          46267 => x"00", -- $0b4bb
          46268 => x"00", -- $0b4bc
          46269 => x"00", -- $0b4bd
          46270 => x"00", -- $0b4be
          46271 => x"00", -- $0b4bf
          46272 => x"00", -- $0b4c0
          46273 => x"00", -- $0b4c1
          46274 => x"00", -- $0b4c2
          46275 => x"00", -- $0b4c3
          46276 => x"00", -- $0b4c4
          46277 => x"00", -- $0b4c5
          46278 => x"00", -- $0b4c6
          46279 => x"00", -- $0b4c7
          46280 => x"00", -- $0b4c8
          46281 => x"00", -- $0b4c9
          46282 => x"00", -- $0b4ca
          46283 => x"00", -- $0b4cb
          46284 => x"00", -- $0b4cc
          46285 => x"00", -- $0b4cd
          46286 => x"00", -- $0b4ce
          46287 => x"00", -- $0b4cf
          46288 => x"00", -- $0b4d0
          46289 => x"00", -- $0b4d1
          46290 => x"00", -- $0b4d2
          46291 => x"00", -- $0b4d3
          46292 => x"00", -- $0b4d4
          46293 => x"00", -- $0b4d5
          46294 => x"00", -- $0b4d6
          46295 => x"00", -- $0b4d7
          46296 => x"00", -- $0b4d8
          46297 => x"00", -- $0b4d9
          46298 => x"00", -- $0b4da
          46299 => x"00", -- $0b4db
          46300 => x"00", -- $0b4dc
          46301 => x"00", -- $0b4dd
          46302 => x"00", -- $0b4de
          46303 => x"00", -- $0b4df
          46304 => x"00", -- $0b4e0
          46305 => x"00", -- $0b4e1
          46306 => x"00", -- $0b4e2
          46307 => x"00", -- $0b4e3
          46308 => x"00", -- $0b4e4
          46309 => x"00", -- $0b4e5
          46310 => x"00", -- $0b4e6
          46311 => x"00", -- $0b4e7
          46312 => x"00", -- $0b4e8
          46313 => x"00", -- $0b4e9
          46314 => x"00", -- $0b4ea
          46315 => x"00", -- $0b4eb
          46316 => x"00", -- $0b4ec
          46317 => x"00", -- $0b4ed
          46318 => x"00", -- $0b4ee
          46319 => x"00", -- $0b4ef
          46320 => x"00", -- $0b4f0
          46321 => x"00", -- $0b4f1
          46322 => x"00", -- $0b4f2
          46323 => x"00", -- $0b4f3
          46324 => x"00", -- $0b4f4
          46325 => x"00", -- $0b4f5
          46326 => x"00", -- $0b4f6
          46327 => x"00", -- $0b4f7
          46328 => x"00", -- $0b4f8
          46329 => x"00", -- $0b4f9
          46330 => x"00", -- $0b4fa
          46331 => x"00", -- $0b4fb
          46332 => x"00", -- $0b4fc
          46333 => x"00", -- $0b4fd
          46334 => x"00", -- $0b4fe
          46335 => x"00", -- $0b4ff
          46336 => x"00", -- $0b500
          46337 => x"00", -- $0b501
          46338 => x"00", -- $0b502
          46339 => x"00", -- $0b503
          46340 => x"00", -- $0b504
          46341 => x"00", -- $0b505
          46342 => x"00", -- $0b506
          46343 => x"00", -- $0b507
          46344 => x"00", -- $0b508
          46345 => x"00", -- $0b509
          46346 => x"00", -- $0b50a
          46347 => x"00", -- $0b50b
          46348 => x"00", -- $0b50c
          46349 => x"00", -- $0b50d
          46350 => x"00", -- $0b50e
          46351 => x"00", -- $0b50f
          46352 => x"00", -- $0b510
          46353 => x"00", -- $0b511
          46354 => x"00", -- $0b512
          46355 => x"00", -- $0b513
          46356 => x"00", -- $0b514
          46357 => x"00", -- $0b515
          46358 => x"00", -- $0b516
          46359 => x"00", -- $0b517
          46360 => x"00", -- $0b518
          46361 => x"00", -- $0b519
          46362 => x"00", -- $0b51a
          46363 => x"00", -- $0b51b
          46364 => x"00", -- $0b51c
          46365 => x"00", -- $0b51d
          46366 => x"00", -- $0b51e
          46367 => x"00", -- $0b51f
          46368 => x"00", -- $0b520
          46369 => x"00", -- $0b521
          46370 => x"00", -- $0b522
          46371 => x"00", -- $0b523
          46372 => x"00", -- $0b524
          46373 => x"00", -- $0b525
          46374 => x"00", -- $0b526
          46375 => x"00", -- $0b527
          46376 => x"00", -- $0b528
          46377 => x"00", -- $0b529
          46378 => x"00", -- $0b52a
          46379 => x"00", -- $0b52b
          46380 => x"00", -- $0b52c
          46381 => x"00", -- $0b52d
          46382 => x"00", -- $0b52e
          46383 => x"00", -- $0b52f
          46384 => x"00", -- $0b530
          46385 => x"00", -- $0b531
          46386 => x"00", -- $0b532
          46387 => x"00", -- $0b533
          46388 => x"00", -- $0b534
          46389 => x"00", -- $0b535
          46390 => x"00", -- $0b536
          46391 => x"00", -- $0b537
          46392 => x"00", -- $0b538
          46393 => x"00", -- $0b539
          46394 => x"00", -- $0b53a
          46395 => x"00", -- $0b53b
          46396 => x"00", -- $0b53c
          46397 => x"00", -- $0b53d
          46398 => x"00", -- $0b53e
          46399 => x"00", -- $0b53f
          46400 => x"00", -- $0b540
          46401 => x"00", -- $0b541
          46402 => x"00", -- $0b542
          46403 => x"00", -- $0b543
          46404 => x"00", -- $0b544
          46405 => x"00", -- $0b545
          46406 => x"00", -- $0b546
          46407 => x"00", -- $0b547
          46408 => x"00", -- $0b548
          46409 => x"00", -- $0b549
          46410 => x"00", -- $0b54a
          46411 => x"00", -- $0b54b
          46412 => x"00", -- $0b54c
          46413 => x"00", -- $0b54d
          46414 => x"00", -- $0b54e
          46415 => x"00", -- $0b54f
          46416 => x"00", -- $0b550
          46417 => x"00", -- $0b551
          46418 => x"00", -- $0b552
          46419 => x"00", -- $0b553
          46420 => x"00", -- $0b554
          46421 => x"00", -- $0b555
          46422 => x"00", -- $0b556
          46423 => x"00", -- $0b557
          46424 => x"00", -- $0b558
          46425 => x"00", -- $0b559
          46426 => x"00", -- $0b55a
          46427 => x"00", -- $0b55b
          46428 => x"00", -- $0b55c
          46429 => x"00", -- $0b55d
          46430 => x"00", -- $0b55e
          46431 => x"00", -- $0b55f
          46432 => x"00", -- $0b560
          46433 => x"00", -- $0b561
          46434 => x"00", -- $0b562
          46435 => x"00", -- $0b563
          46436 => x"00", -- $0b564
          46437 => x"00", -- $0b565
          46438 => x"00", -- $0b566
          46439 => x"00", -- $0b567
          46440 => x"00", -- $0b568
          46441 => x"00", -- $0b569
          46442 => x"00", -- $0b56a
          46443 => x"00", -- $0b56b
          46444 => x"00", -- $0b56c
          46445 => x"00", -- $0b56d
          46446 => x"00", -- $0b56e
          46447 => x"00", -- $0b56f
          46448 => x"00", -- $0b570
          46449 => x"00", -- $0b571
          46450 => x"00", -- $0b572
          46451 => x"00", -- $0b573
          46452 => x"00", -- $0b574
          46453 => x"00", -- $0b575
          46454 => x"00", -- $0b576
          46455 => x"00", -- $0b577
          46456 => x"00", -- $0b578
          46457 => x"00", -- $0b579
          46458 => x"00", -- $0b57a
          46459 => x"00", -- $0b57b
          46460 => x"00", -- $0b57c
          46461 => x"00", -- $0b57d
          46462 => x"00", -- $0b57e
          46463 => x"00", -- $0b57f
          46464 => x"00", -- $0b580
          46465 => x"00", -- $0b581
          46466 => x"00", -- $0b582
          46467 => x"00", -- $0b583
          46468 => x"00", -- $0b584
          46469 => x"00", -- $0b585
          46470 => x"00", -- $0b586
          46471 => x"00", -- $0b587
          46472 => x"00", -- $0b588
          46473 => x"00", -- $0b589
          46474 => x"00", -- $0b58a
          46475 => x"00", -- $0b58b
          46476 => x"00", -- $0b58c
          46477 => x"00", -- $0b58d
          46478 => x"00", -- $0b58e
          46479 => x"00", -- $0b58f
          46480 => x"00", -- $0b590
          46481 => x"00", -- $0b591
          46482 => x"00", -- $0b592
          46483 => x"00", -- $0b593
          46484 => x"00", -- $0b594
          46485 => x"00", -- $0b595
          46486 => x"00", -- $0b596
          46487 => x"00", -- $0b597
          46488 => x"00", -- $0b598
          46489 => x"00", -- $0b599
          46490 => x"00", -- $0b59a
          46491 => x"00", -- $0b59b
          46492 => x"00", -- $0b59c
          46493 => x"00", -- $0b59d
          46494 => x"00", -- $0b59e
          46495 => x"00", -- $0b59f
          46496 => x"00", -- $0b5a0
          46497 => x"00", -- $0b5a1
          46498 => x"00", -- $0b5a2
          46499 => x"00", -- $0b5a3
          46500 => x"00", -- $0b5a4
          46501 => x"00", -- $0b5a5
          46502 => x"00", -- $0b5a6
          46503 => x"00", -- $0b5a7
          46504 => x"00", -- $0b5a8
          46505 => x"00", -- $0b5a9
          46506 => x"00", -- $0b5aa
          46507 => x"00", -- $0b5ab
          46508 => x"00", -- $0b5ac
          46509 => x"00", -- $0b5ad
          46510 => x"00", -- $0b5ae
          46511 => x"00", -- $0b5af
          46512 => x"00", -- $0b5b0
          46513 => x"00", -- $0b5b1
          46514 => x"00", -- $0b5b2
          46515 => x"00", -- $0b5b3
          46516 => x"00", -- $0b5b4
          46517 => x"00", -- $0b5b5
          46518 => x"00", -- $0b5b6
          46519 => x"00", -- $0b5b7
          46520 => x"00", -- $0b5b8
          46521 => x"00", -- $0b5b9
          46522 => x"00", -- $0b5ba
          46523 => x"00", -- $0b5bb
          46524 => x"00", -- $0b5bc
          46525 => x"00", -- $0b5bd
          46526 => x"00", -- $0b5be
          46527 => x"00", -- $0b5bf
          46528 => x"00", -- $0b5c0
          46529 => x"00", -- $0b5c1
          46530 => x"00", -- $0b5c2
          46531 => x"00", -- $0b5c3
          46532 => x"00", -- $0b5c4
          46533 => x"00", -- $0b5c5
          46534 => x"00", -- $0b5c6
          46535 => x"00", -- $0b5c7
          46536 => x"00", -- $0b5c8
          46537 => x"00", -- $0b5c9
          46538 => x"00", -- $0b5ca
          46539 => x"00", -- $0b5cb
          46540 => x"00", -- $0b5cc
          46541 => x"00", -- $0b5cd
          46542 => x"00", -- $0b5ce
          46543 => x"00", -- $0b5cf
          46544 => x"00", -- $0b5d0
          46545 => x"00", -- $0b5d1
          46546 => x"00", -- $0b5d2
          46547 => x"00", -- $0b5d3
          46548 => x"00", -- $0b5d4
          46549 => x"00", -- $0b5d5
          46550 => x"00", -- $0b5d6
          46551 => x"00", -- $0b5d7
          46552 => x"00", -- $0b5d8
          46553 => x"00", -- $0b5d9
          46554 => x"00", -- $0b5da
          46555 => x"00", -- $0b5db
          46556 => x"00", -- $0b5dc
          46557 => x"00", -- $0b5dd
          46558 => x"00", -- $0b5de
          46559 => x"00", -- $0b5df
          46560 => x"00", -- $0b5e0
          46561 => x"00", -- $0b5e1
          46562 => x"00", -- $0b5e2
          46563 => x"00", -- $0b5e3
          46564 => x"00", -- $0b5e4
          46565 => x"00", -- $0b5e5
          46566 => x"00", -- $0b5e6
          46567 => x"00", -- $0b5e7
          46568 => x"00", -- $0b5e8
          46569 => x"00", -- $0b5e9
          46570 => x"00", -- $0b5ea
          46571 => x"00", -- $0b5eb
          46572 => x"00", -- $0b5ec
          46573 => x"00", -- $0b5ed
          46574 => x"00", -- $0b5ee
          46575 => x"00", -- $0b5ef
          46576 => x"00", -- $0b5f0
          46577 => x"00", -- $0b5f1
          46578 => x"00", -- $0b5f2
          46579 => x"00", -- $0b5f3
          46580 => x"00", -- $0b5f4
          46581 => x"00", -- $0b5f5
          46582 => x"00", -- $0b5f6
          46583 => x"00", -- $0b5f7
          46584 => x"00", -- $0b5f8
          46585 => x"00", -- $0b5f9
          46586 => x"00", -- $0b5fa
          46587 => x"00", -- $0b5fb
          46588 => x"00", -- $0b5fc
          46589 => x"00", -- $0b5fd
          46590 => x"00", -- $0b5fe
          46591 => x"00", -- $0b5ff
          46592 => x"00", -- $0b600
          46593 => x"00", -- $0b601
          46594 => x"00", -- $0b602
          46595 => x"00", -- $0b603
          46596 => x"00", -- $0b604
          46597 => x"00", -- $0b605
          46598 => x"00", -- $0b606
          46599 => x"00", -- $0b607
          46600 => x"00", -- $0b608
          46601 => x"00", -- $0b609
          46602 => x"00", -- $0b60a
          46603 => x"00", -- $0b60b
          46604 => x"00", -- $0b60c
          46605 => x"00", -- $0b60d
          46606 => x"00", -- $0b60e
          46607 => x"00", -- $0b60f
          46608 => x"00", -- $0b610
          46609 => x"00", -- $0b611
          46610 => x"00", -- $0b612
          46611 => x"00", -- $0b613
          46612 => x"00", -- $0b614
          46613 => x"00", -- $0b615
          46614 => x"00", -- $0b616
          46615 => x"00", -- $0b617
          46616 => x"00", -- $0b618
          46617 => x"00", -- $0b619
          46618 => x"00", -- $0b61a
          46619 => x"00", -- $0b61b
          46620 => x"00", -- $0b61c
          46621 => x"00", -- $0b61d
          46622 => x"00", -- $0b61e
          46623 => x"00", -- $0b61f
          46624 => x"00", -- $0b620
          46625 => x"00", -- $0b621
          46626 => x"00", -- $0b622
          46627 => x"00", -- $0b623
          46628 => x"00", -- $0b624
          46629 => x"00", -- $0b625
          46630 => x"00", -- $0b626
          46631 => x"00", -- $0b627
          46632 => x"00", -- $0b628
          46633 => x"00", -- $0b629
          46634 => x"00", -- $0b62a
          46635 => x"00", -- $0b62b
          46636 => x"00", -- $0b62c
          46637 => x"00", -- $0b62d
          46638 => x"00", -- $0b62e
          46639 => x"00", -- $0b62f
          46640 => x"00", -- $0b630
          46641 => x"00", -- $0b631
          46642 => x"00", -- $0b632
          46643 => x"00", -- $0b633
          46644 => x"00", -- $0b634
          46645 => x"00", -- $0b635
          46646 => x"00", -- $0b636
          46647 => x"00", -- $0b637
          46648 => x"00", -- $0b638
          46649 => x"00", -- $0b639
          46650 => x"00", -- $0b63a
          46651 => x"00", -- $0b63b
          46652 => x"00", -- $0b63c
          46653 => x"00", -- $0b63d
          46654 => x"00", -- $0b63e
          46655 => x"00", -- $0b63f
          46656 => x"00", -- $0b640
          46657 => x"00", -- $0b641
          46658 => x"00", -- $0b642
          46659 => x"00", -- $0b643
          46660 => x"00", -- $0b644
          46661 => x"00", -- $0b645
          46662 => x"00", -- $0b646
          46663 => x"00", -- $0b647
          46664 => x"00", -- $0b648
          46665 => x"00", -- $0b649
          46666 => x"00", -- $0b64a
          46667 => x"00", -- $0b64b
          46668 => x"00", -- $0b64c
          46669 => x"00", -- $0b64d
          46670 => x"00", -- $0b64e
          46671 => x"00", -- $0b64f
          46672 => x"00", -- $0b650
          46673 => x"00", -- $0b651
          46674 => x"00", -- $0b652
          46675 => x"00", -- $0b653
          46676 => x"00", -- $0b654
          46677 => x"00", -- $0b655
          46678 => x"00", -- $0b656
          46679 => x"00", -- $0b657
          46680 => x"00", -- $0b658
          46681 => x"00", -- $0b659
          46682 => x"00", -- $0b65a
          46683 => x"00", -- $0b65b
          46684 => x"00", -- $0b65c
          46685 => x"00", -- $0b65d
          46686 => x"00", -- $0b65e
          46687 => x"00", -- $0b65f
          46688 => x"00", -- $0b660
          46689 => x"00", -- $0b661
          46690 => x"00", -- $0b662
          46691 => x"00", -- $0b663
          46692 => x"00", -- $0b664
          46693 => x"00", -- $0b665
          46694 => x"00", -- $0b666
          46695 => x"00", -- $0b667
          46696 => x"00", -- $0b668
          46697 => x"00", -- $0b669
          46698 => x"00", -- $0b66a
          46699 => x"00", -- $0b66b
          46700 => x"00", -- $0b66c
          46701 => x"00", -- $0b66d
          46702 => x"00", -- $0b66e
          46703 => x"00", -- $0b66f
          46704 => x"00", -- $0b670
          46705 => x"00", -- $0b671
          46706 => x"00", -- $0b672
          46707 => x"00", -- $0b673
          46708 => x"00", -- $0b674
          46709 => x"00", -- $0b675
          46710 => x"00", -- $0b676
          46711 => x"00", -- $0b677
          46712 => x"00", -- $0b678
          46713 => x"00", -- $0b679
          46714 => x"00", -- $0b67a
          46715 => x"00", -- $0b67b
          46716 => x"00", -- $0b67c
          46717 => x"00", -- $0b67d
          46718 => x"00", -- $0b67e
          46719 => x"00", -- $0b67f
          46720 => x"00", -- $0b680
          46721 => x"00", -- $0b681
          46722 => x"00", -- $0b682
          46723 => x"00", -- $0b683
          46724 => x"00", -- $0b684
          46725 => x"00", -- $0b685
          46726 => x"00", -- $0b686
          46727 => x"00", -- $0b687
          46728 => x"00", -- $0b688
          46729 => x"00", -- $0b689
          46730 => x"00", -- $0b68a
          46731 => x"00", -- $0b68b
          46732 => x"00", -- $0b68c
          46733 => x"00", -- $0b68d
          46734 => x"00", -- $0b68e
          46735 => x"00", -- $0b68f
          46736 => x"00", -- $0b690
          46737 => x"00", -- $0b691
          46738 => x"00", -- $0b692
          46739 => x"00", -- $0b693
          46740 => x"00", -- $0b694
          46741 => x"00", -- $0b695
          46742 => x"00", -- $0b696
          46743 => x"00", -- $0b697
          46744 => x"00", -- $0b698
          46745 => x"00", -- $0b699
          46746 => x"00", -- $0b69a
          46747 => x"00", -- $0b69b
          46748 => x"00", -- $0b69c
          46749 => x"00", -- $0b69d
          46750 => x"00", -- $0b69e
          46751 => x"00", -- $0b69f
          46752 => x"00", -- $0b6a0
          46753 => x"00", -- $0b6a1
          46754 => x"00", -- $0b6a2
          46755 => x"00", -- $0b6a3
          46756 => x"00", -- $0b6a4
          46757 => x"00", -- $0b6a5
          46758 => x"00", -- $0b6a6
          46759 => x"00", -- $0b6a7
          46760 => x"00", -- $0b6a8
          46761 => x"00", -- $0b6a9
          46762 => x"00", -- $0b6aa
          46763 => x"00", -- $0b6ab
          46764 => x"00", -- $0b6ac
          46765 => x"00", -- $0b6ad
          46766 => x"00", -- $0b6ae
          46767 => x"00", -- $0b6af
          46768 => x"00", -- $0b6b0
          46769 => x"00", -- $0b6b1
          46770 => x"00", -- $0b6b2
          46771 => x"00", -- $0b6b3
          46772 => x"00", -- $0b6b4
          46773 => x"00", -- $0b6b5
          46774 => x"00", -- $0b6b6
          46775 => x"00", -- $0b6b7
          46776 => x"00", -- $0b6b8
          46777 => x"00", -- $0b6b9
          46778 => x"00", -- $0b6ba
          46779 => x"00", -- $0b6bb
          46780 => x"00", -- $0b6bc
          46781 => x"00", -- $0b6bd
          46782 => x"00", -- $0b6be
          46783 => x"00", -- $0b6bf
          46784 => x"00", -- $0b6c0
          46785 => x"00", -- $0b6c1
          46786 => x"00", -- $0b6c2
          46787 => x"00", -- $0b6c3
          46788 => x"00", -- $0b6c4
          46789 => x"00", -- $0b6c5
          46790 => x"00", -- $0b6c6
          46791 => x"00", -- $0b6c7
          46792 => x"00", -- $0b6c8
          46793 => x"00", -- $0b6c9
          46794 => x"00", -- $0b6ca
          46795 => x"00", -- $0b6cb
          46796 => x"00", -- $0b6cc
          46797 => x"00", -- $0b6cd
          46798 => x"00", -- $0b6ce
          46799 => x"00", -- $0b6cf
          46800 => x"00", -- $0b6d0
          46801 => x"00", -- $0b6d1
          46802 => x"00", -- $0b6d2
          46803 => x"00", -- $0b6d3
          46804 => x"00", -- $0b6d4
          46805 => x"00", -- $0b6d5
          46806 => x"00", -- $0b6d6
          46807 => x"00", -- $0b6d7
          46808 => x"00", -- $0b6d8
          46809 => x"00", -- $0b6d9
          46810 => x"00", -- $0b6da
          46811 => x"00", -- $0b6db
          46812 => x"00", -- $0b6dc
          46813 => x"00", -- $0b6dd
          46814 => x"00", -- $0b6de
          46815 => x"00", -- $0b6df
          46816 => x"00", -- $0b6e0
          46817 => x"00", -- $0b6e1
          46818 => x"00", -- $0b6e2
          46819 => x"00", -- $0b6e3
          46820 => x"00", -- $0b6e4
          46821 => x"00", -- $0b6e5
          46822 => x"00", -- $0b6e6
          46823 => x"00", -- $0b6e7
          46824 => x"00", -- $0b6e8
          46825 => x"00", -- $0b6e9
          46826 => x"00", -- $0b6ea
          46827 => x"00", -- $0b6eb
          46828 => x"00", -- $0b6ec
          46829 => x"00", -- $0b6ed
          46830 => x"00", -- $0b6ee
          46831 => x"00", -- $0b6ef
          46832 => x"00", -- $0b6f0
          46833 => x"00", -- $0b6f1
          46834 => x"00", -- $0b6f2
          46835 => x"00", -- $0b6f3
          46836 => x"00", -- $0b6f4
          46837 => x"00", -- $0b6f5
          46838 => x"00", -- $0b6f6
          46839 => x"00", -- $0b6f7
          46840 => x"00", -- $0b6f8
          46841 => x"00", -- $0b6f9
          46842 => x"00", -- $0b6fa
          46843 => x"00", -- $0b6fb
          46844 => x"00", -- $0b6fc
          46845 => x"00", -- $0b6fd
          46846 => x"00", -- $0b6fe
          46847 => x"00", -- $0b6ff
          46848 => x"00", -- $0b700
          46849 => x"00", -- $0b701
          46850 => x"00", -- $0b702
          46851 => x"00", -- $0b703
          46852 => x"00", -- $0b704
          46853 => x"00", -- $0b705
          46854 => x"00", -- $0b706
          46855 => x"00", -- $0b707
          46856 => x"00", -- $0b708
          46857 => x"00", -- $0b709
          46858 => x"00", -- $0b70a
          46859 => x"00", -- $0b70b
          46860 => x"00", -- $0b70c
          46861 => x"00", -- $0b70d
          46862 => x"00", -- $0b70e
          46863 => x"00", -- $0b70f
          46864 => x"00", -- $0b710
          46865 => x"00", -- $0b711
          46866 => x"00", -- $0b712
          46867 => x"00", -- $0b713
          46868 => x"00", -- $0b714
          46869 => x"00", -- $0b715
          46870 => x"00", -- $0b716
          46871 => x"00", -- $0b717
          46872 => x"00", -- $0b718
          46873 => x"00", -- $0b719
          46874 => x"00", -- $0b71a
          46875 => x"00", -- $0b71b
          46876 => x"00", -- $0b71c
          46877 => x"00", -- $0b71d
          46878 => x"00", -- $0b71e
          46879 => x"00", -- $0b71f
          46880 => x"00", -- $0b720
          46881 => x"00", -- $0b721
          46882 => x"00", -- $0b722
          46883 => x"00", -- $0b723
          46884 => x"00", -- $0b724
          46885 => x"00", -- $0b725
          46886 => x"00", -- $0b726
          46887 => x"00", -- $0b727
          46888 => x"00", -- $0b728
          46889 => x"00", -- $0b729
          46890 => x"00", -- $0b72a
          46891 => x"00", -- $0b72b
          46892 => x"00", -- $0b72c
          46893 => x"00", -- $0b72d
          46894 => x"00", -- $0b72e
          46895 => x"00", -- $0b72f
          46896 => x"00", -- $0b730
          46897 => x"00", -- $0b731
          46898 => x"00", -- $0b732
          46899 => x"00", -- $0b733
          46900 => x"00", -- $0b734
          46901 => x"00", -- $0b735
          46902 => x"00", -- $0b736
          46903 => x"00", -- $0b737
          46904 => x"00", -- $0b738
          46905 => x"00", -- $0b739
          46906 => x"00", -- $0b73a
          46907 => x"00", -- $0b73b
          46908 => x"00", -- $0b73c
          46909 => x"00", -- $0b73d
          46910 => x"00", -- $0b73e
          46911 => x"00", -- $0b73f
          46912 => x"00", -- $0b740
          46913 => x"00", -- $0b741
          46914 => x"00", -- $0b742
          46915 => x"00", -- $0b743
          46916 => x"00", -- $0b744
          46917 => x"00", -- $0b745
          46918 => x"00", -- $0b746
          46919 => x"00", -- $0b747
          46920 => x"00", -- $0b748
          46921 => x"00", -- $0b749
          46922 => x"00", -- $0b74a
          46923 => x"00", -- $0b74b
          46924 => x"00", -- $0b74c
          46925 => x"00", -- $0b74d
          46926 => x"00", -- $0b74e
          46927 => x"00", -- $0b74f
          46928 => x"00", -- $0b750
          46929 => x"00", -- $0b751
          46930 => x"00", -- $0b752
          46931 => x"00", -- $0b753
          46932 => x"00", -- $0b754
          46933 => x"00", -- $0b755
          46934 => x"00", -- $0b756
          46935 => x"00", -- $0b757
          46936 => x"00", -- $0b758
          46937 => x"00", -- $0b759
          46938 => x"00", -- $0b75a
          46939 => x"00", -- $0b75b
          46940 => x"00", -- $0b75c
          46941 => x"00", -- $0b75d
          46942 => x"00", -- $0b75e
          46943 => x"00", -- $0b75f
          46944 => x"00", -- $0b760
          46945 => x"00", -- $0b761
          46946 => x"00", -- $0b762
          46947 => x"00", -- $0b763
          46948 => x"00", -- $0b764
          46949 => x"00", -- $0b765
          46950 => x"00", -- $0b766
          46951 => x"00", -- $0b767
          46952 => x"00", -- $0b768
          46953 => x"00", -- $0b769
          46954 => x"00", -- $0b76a
          46955 => x"00", -- $0b76b
          46956 => x"00", -- $0b76c
          46957 => x"00", -- $0b76d
          46958 => x"00", -- $0b76e
          46959 => x"00", -- $0b76f
          46960 => x"00", -- $0b770
          46961 => x"00", -- $0b771
          46962 => x"00", -- $0b772
          46963 => x"00", -- $0b773
          46964 => x"00", -- $0b774
          46965 => x"00", -- $0b775
          46966 => x"00", -- $0b776
          46967 => x"00", -- $0b777
          46968 => x"00", -- $0b778
          46969 => x"00", -- $0b779
          46970 => x"00", -- $0b77a
          46971 => x"00", -- $0b77b
          46972 => x"00", -- $0b77c
          46973 => x"00", -- $0b77d
          46974 => x"00", -- $0b77e
          46975 => x"00", -- $0b77f
          46976 => x"00", -- $0b780
          46977 => x"00", -- $0b781
          46978 => x"00", -- $0b782
          46979 => x"00", -- $0b783
          46980 => x"00", -- $0b784
          46981 => x"00", -- $0b785
          46982 => x"00", -- $0b786
          46983 => x"00", -- $0b787
          46984 => x"00", -- $0b788
          46985 => x"00", -- $0b789
          46986 => x"00", -- $0b78a
          46987 => x"00", -- $0b78b
          46988 => x"00", -- $0b78c
          46989 => x"00", -- $0b78d
          46990 => x"00", -- $0b78e
          46991 => x"00", -- $0b78f
          46992 => x"00", -- $0b790
          46993 => x"00", -- $0b791
          46994 => x"00", -- $0b792
          46995 => x"00", -- $0b793
          46996 => x"00", -- $0b794
          46997 => x"00", -- $0b795
          46998 => x"00", -- $0b796
          46999 => x"00", -- $0b797
          47000 => x"00", -- $0b798
          47001 => x"00", -- $0b799
          47002 => x"00", -- $0b79a
          47003 => x"00", -- $0b79b
          47004 => x"00", -- $0b79c
          47005 => x"00", -- $0b79d
          47006 => x"00", -- $0b79e
          47007 => x"00", -- $0b79f
          47008 => x"00", -- $0b7a0
          47009 => x"00", -- $0b7a1
          47010 => x"00", -- $0b7a2
          47011 => x"00", -- $0b7a3
          47012 => x"00", -- $0b7a4
          47013 => x"00", -- $0b7a5
          47014 => x"00", -- $0b7a6
          47015 => x"00", -- $0b7a7
          47016 => x"00", -- $0b7a8
          47017 => x"00", -- $0b7a9
          47018 => x"00", -- $0b7aa
          47019 => x"00", -- $0b7ab
          47020 => x"00", -- $0b7ac
          47021 => x"00", -- $0b7ad
          47022 => x"00", -- $0b7ae
          47023 => x"00", -- $0b7af
          47024 => x"00", -- $0b7b0
          47025 => x"00", -- $0b7b1
          47026 => x"00", -- $0b7b2
          47027 => x"00", -- $0b7b3
          47028 => x"00", -- $0b7b4
          47029 => x"00", -- $0b7b5
          47030 => x"00", -- $0b7b6
          47031 => x"00", -- $0b7b7
          47032 => x"00", -- $0b7b8
          47033 => x"00", -- $0b7b9
          47034 => x"00", -- $0b7ba
          47035 => x"00", -- $0b7bb
          47036 => x"00", -- $0b7bc
          47037 => x"00", -- $0b7bd
          47038 => x"00", -- $0b7be
          47039 => x"00", -- $0b7bf
          47040 => x"00", -- $0b7c0
          47041 => x"00", -- $0b7c1
          47042 => x"00", -- $0b7c2
          47043 => x"00", -- $0b7c3
          47044 => x"00", -- $0b7c4
          47045 => x"00", -- $0b7c5
          47046 => x"00", -- $0b7c6
          47047 => x"00", -- $0b7c7
          47048 => x"00", -- $0b7c8
          47049 => x"00", -- $0b7c9
          47050 => x"00", -- $0b7ca
          47051 => x"00", -- $0b7cb
          47052 => x"00", -- $0b7cc
          47053 => x"00", -- $0b7cd
          47054 => x"00", -- $0b7ce
          47055 => x"00", -- $0b7cf
          47056 => x"00", -- $0b7d0
          47057 => x"00", -- $0b7d1
          47058 => x"00", -- $0b7d2
          47059 => x"00", -- $0b7d3
          47060 => x"00", -- $0b7d4
          47061 => x"00", -- $0b7d5
          47062 => x"00", -- $0b7d6
          47063 => x"00", -- $0b7d7
          47064 => x"00", -- $0b7d8
          47065 => x"00", -- $0b7d9
          47066 => x"00", -- $0b7da
          47067 => x"00", -- $0b7db
          47068 => x"00", -- $0b7dc
          47069 => x"00", -- $0b7dd
          47070 => x"00", -- $0b7de
          47071 => x"00", -- $0b7df
          47072 => x"00", -- $0b7e0
          47073 => x"00", -- $0b7e1
          47074 => x"00", -- $0b7e2
          47075 => x"00", -- $0b7e3
          47076 => x"00", -- $0b7e4
          47077 => x"00", -- $0b7e5
          47078 => x"00", -- $0b7e6
          47079 => x"00", -- $0b7e7
          47080 => x"00", -- $0b7e8
          47081 => x"00", -- $0b7e9
          47082 => x"00", -- $0b7ea
          47083 => x"00", -- $0b7eb
          47084 => x"00", -- $0b7ec
          47085 => x"00", -- $0b7ed
          47086 => x"00", -- $0b7ee
          47087 => x"00", -- $0b7ef
          47088 => x"00", -- $0b7f0
          47089 => x"00", -- $0b7f1
          47090 => x"00", -- $0b7f2
          47091 => x"00", -- $0b7f3
          47092 => x"00", -- $0b7f4
          47093 => x"00", -- $0b7f5
          47094 => x"00", -- $0b7f6
          47095 => x"00", -- $0b7f7
          47096 => x"00", -- $0b7f8
          47097 => x"00", -- $0b7f9
          47098 => x"00", -- $0b7fa
          47099 => x"00", -- $0b7fb
          47100 => x"00", -- $0b7fc
          47101 => x"00", -- $0b7fd
          47102 => x"00", -- $0b7fe
          47103 => x"00", -- $0b7ff
          47104 => x"00", -- $0b800
          47105 => x"00", -- $0b801
          47106 => x"00", -- $0b802
          47107 => x"00", -- $0b803
          47108 => x"00", -- $0b804
          47109 => x"00", -- $0b805
          47110 => x"00", -- $0b806
          47111 => x"00", -- $0b807
          47112 => x"00", -- $0b808
          47113 => x"00", -- $0b809
          47114 => x"00", -- $0b80a
          47115 => x"00", -- $0b80b
          47116 => x"00", -- $0b80c
          47117 => x"00", -- $0b80d
          47118 => x"00", -- $0b80e
          47119 => x"00", -- $0b80f
          47120 => x"00", -- $0b810
          47121 => x"00", -- $0b811
          47122 => x"00", -- $0b812
          47123 => x"00", -- $0b813
          47124 => x"00", -- $0b814
          47125 => x"00", -- $0b815
          47126 => x"00", -- $0b816
          47127 => x"00", -- $0b817
          47128 => x"00", -- $0b818
          47129 => x"00", -- $0b819
          47130 => x"00", -- $0b81a
          47131 => x"00", -- $0b81b
          47132 => x"00", -- $0b81c
          47133 => x"00", -- $0b81d
          47134 => x"00", -- $0b81e
          47135 => x"00", -- $0b81f
          47136 => x"00", -- $0b820
          47137 => x"00", -- $0b821
          47138 => x"00", -- $0b822
          47139 => x"00", -- $0b823
          47140 => x"00", -- $0b824
          47141 => x"00", -- $0b825
          47142 => x"00", -- $0b826
          47143 => x"00", -- $0b827
          47144 => x"00", -- $0b828
          47145 => x"00", -- $0b829
          47146 => x"00", -- $0b82a
          47147 => x"00", -- $0b82b
          47148 => x"00", -- $0b82c
          47149 => x"00", -- $0b82d
          47150 => x"00", -- $0b82e
          47151 => x"00", -- $0b82f
          47152 => x"00", -- $0b830
          47153 => x"00", -- $0b831
          47154 => x"00", -- $0b832
          47155 => x"00", -- $0b833
          47156 => x"00", -- $0b834
          47157 => x"00", -- $0b835
          47158 => x"00", -- $0b836
          47159 => x"00", -- $0b837
          47160 => x"00", -- $0b838
          47161 => x"00", -- $0b839
          47162 => x"00", -- $0b83a
          47163 => x"00", -- $0b83b
          47164 => x"00", -- $0b83c
          47165 => x"00", -- $0b83d
          47166 => x"00", -- $0b83e
          47167 => x"00", -- $0b83f
          47168 => x"00", -- $0b840
          47169 => x"00", -- $0b841
          47170 => x"00", -- $0b842
          47171 => x"00", -- $0b843
          47172 => x"00", -- $0b844
          47173 => x"00", -- $0b845
          47174 => x"00", -- $0b846
          47175 => x"00", -- $0b847
          47176 => x"00", -- $0b848
          47177 => x"00", -- $0b849
          47178 => x"00", -- $0b84a
          47179 => x"00", -- $0b84b
          47180 => x"00", -- $0b84c
          47181 => x"00", -- $0b84d
          47182 => x"00", -- $0b84e
          47183 => x"00", -- $0b84f
          47184 => x"00", -- $0b850
          47185 => x"00", -- $0b851
          47186 => x"00", -- $0b852
          47187 => x"00", -- $0b853
          47188 => x"00", -- $0b854
          47189 => x"00", -- $0b855
          47190 => x"00", -- $0b856
          47191 => x"00", -- $0b857
          47192 => x"00", -- $0b858
          47193 => x"00", -- $0b859
          47194 => x"00", -- $0b85a
          47195 => x"00", -- $0b85b
          47196 => x"00", -- $0b85c
          47197 => x"00", -- $0b85d
          47198 => x"00", -- $0b85e
          47199 => x"00", -- $0b85f
          47200 => x"00", -- $0b860
          47201 => x"00", -- $0b861
          47202 => x"00", -- $0b862
          47203 => x"00", -- $0b863
          47204 => x"00", -- $0b864
          47205 => x"00", -- $0b865
          47206 => x"00", -- $0b866
          47207 => x"00", -- $0b867
          47208 => x"00", -- $0b868
          47209 => x"00", -- $0b869
          47210 => x"00", -- $0b86a
          47211 => x"00", -- $0b86b
          47212 => x"00", -- $0b86c
          47213 => x"00", -- $0b86d
          47214 => x"00", -- $0b86e
          47215 => x"00", -- $0b86f
          47216 => x"00", -- $0b870
          47217 => x"00", -- $0b871
          47218 => x"00", -- $0b872
          47219 => x"00", -- $0b873
          47220 => x"00", -- $0b874
          47221 => x"00", -- $0b875
          47222 => x"00", -- $0b876
          47223 => x"00", -- $0b877
          47224 => x"00", -- $0b878
          47225 => x"00", -- $0b879
          47226 => x"00", -- $0b87a
          47227 => x"00", -- $0b87b
          47228 => x"00", -- $0b87c
          47229 => x"00", -- $0b87d
          47230 => x"00", -- $0b87e
          47231 => x"00", -- $0b87f
          47232 => x"00", -- $0b880
          47233 => x"00", -- $0b881
          47234 => x"00", -- $0b882
          47235 => x"00", -- $0b883
          47236 => x"00", -- $0b884
          47237 => x"00", -- $0b885
          47238 => x"00", -- $0b886
          47239 => x"00", -- $0b887
          47240 => x"00", -- $0b888
          47241 => x"00", -- $0b889
          47242 => x"00", -- $0b88a
          47243 => x"00", -- $0b88b
          47244 => x"00", -- $0b88c
          47245 => x"00", -- $0b88d
          47246 => x"00", -- $0b88e
          47247 => x"00", -- $0b88f
          47248 => x"00", -- $0b890
          47249 => x"00", -- $0b891
          47250 => x"00", -- $0b892
          47251 => x"00", -- $0b893
          47252 => x"00", -- $0b894
          47253 => x"00", -- $0b895
          47254 => x"00", -- $0b896
          47255 => x"00", -- $0b897
          47256 => x"00", -- $0b898
          47257 => x"00", -- $0b899
          47258 => x"00", -- $0b89a
          47259 => x"00", -- $0b89b
          47260 => x"00", -- $0b89c
          47261 => x"00", -- $0b89d
          47262 => x"00", -- $0b89e
          47263 => x"00", -- $0b89f
          47264 => x"00", -- $0b8a0
          47265 => x"00", -- $0b8a1
          47266 => x"00", -- $0b8a2
          47267 => x"00", -- $0b8a3
          47268 => x"00", -- $0b8a4
          47269 => x"00", -- $0b8a5
          47270 => x"00", -- $0b8a6
          47271 => x"00", -- $0b8a7
          47272 => x"00", -- $0b8a8
          47273 => x"00", -- $0b8a9
          47274 => x"00", -- $0b8aa
          47275 => x"00", -- $0b8ab
          47276 => x"00", -- $0b8ac
          47277 => x"00", -- $0b8ad
          47278 => x"00", -- $0b8ae
          47279 => x"00", -- $0b8af
          47280 => x"00", -- $0b8b0
          47281 => x"00", -- $0b8b1
          47282 => x"00", -- $0b8b2
          47283 => x"00", -- $0b8b3
          47284 => x"00", -- $0b8b4
          47285 => x"00", -- $0b8b5
          47286 => x"00", -- $0b8b6
          47287 => x"00", -- $0b8b7
          47288 => x"00", -- $0b8b8
          47289 => x"00", -- $0b8b9
          47290 => x"00", -- $0b8ba
          47291 => x"00", -- $0b8bb
          47292 => x"00", -- $0b8bc
          47293 => x"00", -- $0b8bd
          47294 => x"00", -- $0b8be
          47295 => x"00", -- $0b8bf
          47296 => x"00", -- $0b8c0
          47297 => x"00", -- $0b8c1
          47298 => x"00", -- $0b8c2
          47299 => x"00", -- $0b8c3
          47300 => x"00", -- $0b8c4
          47301 => x"00", -- $0b8c5
          47302 => x"00", -- $0b8c6
          47303 => x"00", -- $0b8c7
          47304 => x"00", -- $0b8c8
          47305 => x"00", -- $0b8c9
          47306 => x"00", -- $0b8ca
          47307 => x"00", -- $0b8cb
          47308 => x"00", -- $0b8cc
          47309 => x"00", -- $0b8cd
          47310 => x"00", -- $0b8ce
          47311 => x"00", -- $0b8cf
          47312 => x"00", -- $0b8d0
          47313 => x"00", -- $0b8d1
          47314 => x"00", -- $0b8d2
          47315 => x"00", -- $0b8d3
          47316 => x"00", -- $0b8d4
          47317 => x"00", -- $0b8d5
          47318 => x"00", -- $0b8d6
          47319 => x"00", -- $0b8d7
          47320 => x"00", -- $0b8d8
          47321 => x"00", -- $0b8d9
          47322 => x"00", -- $0b8da
          47323 => x"00", -- $0b8db
          47324 => x"00", -- $0b8dc
          47325 => x"00", -- $0b8dd
          47326 => x"00", -- $0b8de
          47327 => x"00", -- $0b8df
          47328 => x"00", -- $0b8e0
          47329 => x"00", -- $0b8e1
          47330 => x"00", -- $0b8e2
          47331 => x"00", -- $0b8e3
          47332 => x"00", -- $0b8e4
          47333 => x"00", -- $0b8e5
          47334 => x"00", -- $0b8e6
          47335 => x"00", -- $0b8e7
          47336 => x"00", -- $0b8e8
          47337 => x"00", -- $0b8e9
          47338 => x"00", -- $0b8ea
          47339 => x"00", -- $0b8eb
          47340 => x"00", -- $0b8ec
          47341 => x"00", -- $0b8ed
          47342 => x"00", -- $0b8ee
          47343 => x"00", -- $0b8ef
          47344 => x"00", -- $0b8f0
          47345 => x"00", -- $0b8f1
          47346 => x"00", -- $0b8f2
          47347 => x"00", -- $0b8f3
          47348 => x"00", -- $0b8f4
          47349 => x"00", -- $0b8f5
          47350 => x"00", -- $0b8f6
          47351 => x"00", -- $0b8f7
          47352 => x"00", -- $0b8f8
          47353 => x"00", -- $0b8f9
          47354 => x"00", -- $0b8fa
          47355 => x"00", -- $0b8fb
          47356 => x"00", -- $0b8fc
          47357 => x"00", -- $0b8fd
          47358 => x"00", -- $0b8fe
          47359 => x"00", -- $0b8ff
          47360 => x"00", -- $0b900
          47361 => x"00", -- $0b901
          47362 => x"00", -- $0b902
          47363 => x"00", -- $0b903
          47364 => x"00", -- $0b904
          47365 => x"00", -- $0b905
          47366 => x"00", -- $0b906
          47367 => x"00", -- $0b907
          47368 => x"00", -- $0b908
          47369 => x"00", -- $0b909
          47370 => x"00", -- $0b90a
          47371 => x"00", -- $0b90b
          47372 => x"00", -- $0b90c
          47373 => x"00", -- $0b90d
          47374 => x"00", -- $0b90e
          47375 => x"00", -- $0b90f
          47376 => x"00", -- $0b910
          47377 => x"00", -- $0b911
          47378 => x"00", -- $0b912
          47379 => x"00", -- $0b913
          47380 => x"00", -- $0b914
          47381 => x"00", -- $0b915
          47382 => x"00", -- $0b916
          47383 => x"00", -- $0b917
          47384 => x"00", -- $0b918
          47385 => x"00", -- $0b919
          47386 => x"00", -- $0b91a
          47387 => x"00", -- $0b91b
          47388 => x"00", -- $0b91c
          47389 => x"00", -- $0b91d
          47390 => x"00", -- $0b91e
          47391 => x"00", -- $0b91f
          47392 => x"00", -- $0b920
          47393 => x"00", -- $0b921
          47394 => x"00", -- $0b922
          47395 => x"00", -- $0b923
          47396 => x"00", -- $0b924
          47397 => x"00", -- $0b925
          47398 => x"00", -- $0b926
          47399 => x"00", -- $0b927
          47400 => x"00", -- $0b928
          47401 => x"00", -- $0b929
          47402 => x"00", -- $0b92a
          47403 => x"00", -- $0b92b
          47404 => x"00", -- $0b92c
          47405 => x"00", -- $0b92d
          47406 => x"00", -- $0b92e
          47407 => x"00", -- $0b92f
          47408 => x"00", -- $0b930
          47409 => x"00", -- $0b931
          47410 => x"00", -- $0b932
          47411 => x"00", -- $0b933
          47412 => x"00", -- $0b934
          47413 => x"00", -- $0b935
          47414 => x"00", -- $0b936
          47415 => x"00", -- $0b937
          47416 => x"00", -- $0b938
          47417 => x"00", -- $0b939
          47418 => x"00", -- $0b93a
          47419 => x"00", -- $0b93b
          47420 => x"00", -- $0b93c
          47421 => x"00", -- $0b93d
          47422 => x"00", -- $0b93e
          47423 => x"00", -- $0b93f
          47424 => x"00", -- $0b940
          47425 => x"00", -- $0b941
          47426 => x"00", -- $0b942
          47427 => x"00", -- $0b943
          47428 => x"00", -- $0b944
          47429 => x"00", -- $0b945
          47430 => x"00", -- $0b946
          47431 => x"00", -- $0b947
          47432 => x"00", -- $0b948
          47433 => x"00", -- $0b949
          47434 => x"00", -- $0b94a
          47435 => x"00", -- $0b94b
          47436 => x"00", -- $0b94c
          47437 => x"00", -- $0b94d
          47438 => x"00", -- $0b94e
          47439 => x"00", -- $0b94f
          47440 => x"00", -- $0b950
          47441 => x"00", -- $0b951
          47442 => x"00", -- $0b952
          47443 => x"00", -- $0b953
          47444 => x"00", -- $0b954
          47445 => x"00", -- $0b955
          47446 => x"00", -- $0b956
          47447 => x"00", -- $0b957
          47448 => x"00", -- $0b958
          47449 => x"00", -- $0b959
          47450 => x"00", -- $0b95a
          47451 => x"00", -- $0b95b
          47452 => x"00", -- $0b95c
          47453 => x"00", -- $0b95d
          47454 => x"00", -- $0b95e
          47455 => x"00", -- $0b95f
          47456 => x"00", -- $0b960
          47457 => x"00", -- $0b961
          47458 => x"00", -- $0b962
          47459 => x"00", -- $0b963
          47460 => x"00", -- $0b964
          47461 => x"00", -- $0b965
          47462 => x"00", -- $0b966
          47463 => x"00", -- $0b967
          47464 => x"00", -- $0b968
          47465 => x"00", -- $0b969
          47466 => x"00", -- $0b96a
          47467 => x"00", -- $0b96b
          47468 => x"00", -- $0b96c
          47469 => x"00", -- $0b96d
          47470 => x"00", -- $0b96e
          47471 => x"00", -- $0b96f
          47472 => x"00", -- $0b970
          47473 => x"00", -- $0b971
          47474 => x"00", -- $0b972
          47475 => x"00", -- $0b973
          47476 => x"00", -- $0b974
          47477 => x"00", -- $0b975
          47478 => x"00", -- $0b976
          47479 => x"00", -- $0b977
          47480 => x"00", -- $0b978
          47481 => x"00", -- $0b979
          47482 => x"00", -- $0b97a
          47483 => x"00", -- $0b97b
          47484 => x"00", -- $0b97c
          47485 => x"00", -- $0b97d
          47486 => x"00", -- $0b97e
          47487 => x"00", -- $0b97f
          47488 => x"00", -- $0b980
          47489 => x"00", -- $0b981
          47490 => x"00", -- $0b982
          47491 => x"00", -- $0b983
          47492 => x"00", -- $0b984
          47493 => x"00", -- $0b985
          47494 => x"00", -- $0b986
          47495 => x"00", -- $0b987
          47496 => x"00", -- $0b988
          47497 => x"00", -- $0b989
          47498 => x"00", -- $0b98a
          47499 => x"00", -- $0b98b
          47500 => x"00", -- $0b98c
          47501 => x"00", -- $0b98d
          47502 => x"00", -- $0b98e
          47503 => x"00", -- $0b98f
          47504 => x"00", -- $0b990
          47505 => x"00", -- $0b991
          47506 => x"00", -- $0b992
          47507 => x"00", -- $0b993
          47508 => x"00", -- $0b994
          47509 => x"00", -- $0b995
          47510 => x"00", -- $0b996
          47511 => x"00", -- $0b997
          47512 => x"00", -- $0b998
          47513 => x"00", -- $0b999
          47514 => x"00", -- $0b99a
          47515 => x"00", -- $0b99b
          47516 => x"00", -- $0b99c
          47517 => x"00", -- $0b99d
          47518 => x"00", -- $0b99e
          47519 => x"00", -- $0b99f
          47520 => x"00", -- $0b9a0
          47521 => x"00", -- $0b9a1
          47522 => x"00", -- $0b9a2
          47523 => x"00", -- $0b9a3
          47524 => x"00", -- $0b9a4
          47525 => x"00", -- $0b9a5
          47526 => x"00", -- $0b9a6
          47527 => x"00", -- $0b9a7
          47528 => x"00", -- $0b9a8
          47529 => x"00", -- $0b9a9
          47530 => x"00", -- $0b9aa
          47531 => x"00", -- $0b9ab
          47532 => x"00", -- $0b9ac
          47533 => x"00", -- $0b9ad
          47534 => x"00", -- $0b9ae
          47535 => x"00", -- $0b9af
          47536 => x"00", -- $0b9b0
          47537 => x"00", -- $0b9b1
          47538 => x"00", -- $0b9b2
          47539 => x"00", -- $0b9b3
          47540 => x"00", -- $0b9b4
          47541 => x"00", -- $0b9b5
          47542 => x"00", -- $0b9b6
          47543 => x"00", -- $0b9b7
          47544 => x"00", -- $0b9b8
          47545 => x"00", -- $0b9b9
          47546 => x"00", -- $0b9ba
          47547 => x"00", -- $0b9bb
          47548 => x"00", -- $0b9bc
          47549 => x"00", -- $0b9bd
          47550 => x"00", -- $0b9be
          47551 => x"00", -- $0b9bf
          47552 => x"00", -- $0b9c0
          47553 => x"00", -- $0b9c1
          47554 => x"00", -- $0b9c2
          47555 => x"00", -- $0b9c3
          47556 => x"00", -- $0b9c4
          47557 => x"00", -- $0b9c5
          47558 => x"00", -- $0b9c6
          47559 => x"00", -- $0b9c7
          47560 => x"00", -- $0b9c8
          47561 => x"00", -- $0b9c9
          47562 => x"00", -- $0b9ca
          47563 => x"00", -- $0b9cb
          47564 => x"00", -- $0b9cc
          47565 => x"00", -- $0b9cd
          47566 => x"00", -- $0b9ce
          47567 => x"00", -- $0b9cf
          47568 => x"00", -- $0b9d0
          47569 => x"00", -- $0b9d1
          47570 => x"00", -- $0b9d2
          47571 => x"00", -- $0b9d3
          47572 => x"00", -- $0b9d4
          47573 => x"00", -- $0b9d5
          47574 => x"00", -- $0b9d6
          47575 => x"00", -- $0b9d7
          47576 => x"00", -- $0b9d8
          47577 => x"00", -- $0b9d9
          47578 => x"00", -- $0b9da
          47579 => x"00", -- $0b9db
          47580 => x"00", -- $0b9dc
          47581 => x"00", -- $0b9dd
          47582 => x"00", -- $0b9de
          47583 => x"00", -- $0b9df
          47584 => x"00", -- $0b9e0
          47585 => x"00", -- $0b9e1
          47586 => x"00", -- $0b9e2
          47587 => x"00", -- $0b9e3
          47588 => x"00", -- $0b9e4
          47589 => x"00", -- $0b9e5
          47590 => x"00", -- $0b9e6
          47591 => x"00", -- $0b9e7
          47592 => x"00", -- $0b9e8
          47593 => x"00", -- $0b9e9
          47594 => x"00", -- $0b9ea
          47595 => x"00", -- $0b9eb
          47596 => x"00", -- $0b9ec
          47597 => x"00", -- $0b9ed
          47598 => x"00", -- $0b9ee
          47599 => x"00", -- $0b9ef
          47600 => x"00", -- $0b9f0
          47601 => x"00", -- $0b9f1
          47602 => x"00", -- $0b9f2
          47603 => x"00", -- $0b9f3
          47604 => x"00", -- $0b9f4
          47605 => x"00", -- $0b9f5
          47606 => x"00", -- $0b9f6
          47607 => x"00", -- $0b9f7
          47608 => x"00", -- $0b9f8
          47609 => x"00", -- $0b9f9
          47610 => x"00", -- $0b9fa
          47611 => x"00", -- $0b9fb
          47612 => x"00", -- $0b9fc
          47613 => x"00", -- $0b9fd
          47614 => x"00", -- $0b9fe
          47615 => x"00", -- $0b9ff
          47616 => x"00", -- $0ba00
          47617 => x"00", -- $0ba01
          47618 => x"00", -- $0ba02
          47619 => x"00", -- $0ba03
          47620 => x"00", -- $0ba04
          47621 => x"00", -- $0ba05
          47622 => x"00", -- $0ba06
          47623 => x"00", -- $0ba07
          47624 => x"00", -- $0ba08
          47625 => x"00", -- $0ba09
          47626 => x"00", -- $0ba0a
          47627 => x"00", -- $0ba0b
          47628 => x"00", -- $0ba0c
          47629 => x"00", -- $0ba0d
          47630 => x"00", -- $0ba0e
          47631 => x"00", -- $0ba0f
          47632 => x"00", -- $0ba10
          47633 => x"00", -- $0ba11
          47634 => x"00", -- $0ba12
          47635 => x"00", -- $0ba13
          47636 => x"00", -- $0ba14
          47637 => x"00", -- $0ba15
          47638 => x"00", -- $0ba16
          47639 => x"00", -- $0ba17
          47640 => x"00", -- $0ba18
          47641 => x"00", -- $0ba19
          47642 => x"00", -- $0ba1a
          47643 => x"00", -- $0ba1b
          47644 => x"00", -- $0ba1c
          47645 => x"00", -- $0ba1d
          47646 => x"00", -- $0ba1e
          47647 => x"00", -- $0ba1f
          47648 => x"00", -- $0ba20
          47649 => x"00", -- $0ba21
          47650 => x"00", -- $0ba22
          47651 => x"00", -- $0ba23
          47652 => x"00", -- $0ba24
          47653 => x"00", -- $0ba25
          47654 => x"00", -- $0ba26
          47655 => x"00", -- $0ba27
          47656 => x"00", -- $0ba28
          47657 => x"00", -- $0ba29
          47658 => x"00", -- $0ba2a
          47659 => x"00", -- $0ba2b
          47660 => x"00", -- $0ba2c
          47661 => x"00", -- $0ba2d
          47662 => x"00", -- $0ba2e
          47663 => x"00", -- $0ba2f
          47664 => x"00", -- $0ba30
          47665 => x"00", -- $0ba31
          47666 => x"00", -- $0ba32
          47667 => x"00", -- $0ba33
          47668 => x"00", -- $0ba34
          47669 => x"00", -- $0ba35
          47670 => x"00", -- $0ba36
          47671 => x"00", -- $0ba37
          47672 => x"00", -- $0ba38
          47673 => x"00", -- $0ba39
          47674 => x"00", -- $0ba3a
          47675 => x"00", -- $0ba3b
          47676 => x"00", -- $0ba3c
          47677 => x"00", -- $0ba3d
          47678 => x"00", -- $0ba3e
          47679 => x"00", -- $0ba3f
          47680 => x"00", -- $0ba40
          47681 => x"00", -- $0ba41
          47682 => x"00", -- $0ba42
          47683 => x"00", -- $0ba43
          47684 => x"00", -- $0ba44
          47685 => x"00", -- $0ba45
          47686 => x"00", -- $0ba46
          47687 => x"00", -- $0ba47
          47688 => x"00", -- $0ba48
          47689 => x"00", -- $0ba49
          47690 => x"00", -- $0ba4a
          47691 => x"00", -- $0ba4b
          47692 => x"00", -- $0ba4c
          47693 => x"00", -- $0ba4d
          47694 => x"00", -- $0ba4e
          47695 => x"00", -- $0ba4f
          47696 => x"00", -- $0ba50
          47697 => x"00", -- $0ba51
          47698 => x"00", -- $0ba52
          47699 => x"00", -- $0ba53
          47700 => x"00", -- $0ba54
          47701 => x"00", -- $0ba55
          47702 => x"00", -- $0ba56
          47703 => x"00", -- $0ba57
          47704 => x"00", -- $0ba58
          47705 => x"00", -- $0ba59
          47706 => x"00", -- $0ba5a
          47707 => x"00", -- $0ba5b
          47708 => x"00", -- $0ba5c
          47709 => x"00", -- $0ba5d
          47710 => x"00", -- $0ba5e
          47711 => x"00", -- $0ba5f
          47712 => x"00", -- $0ba60
          47713 => x"00", -- $0ba61
          47714 => x"00", -- $0ba62
          47715 => x"00", -- $0ba63
          47716 => x"00", -- $0ba64
          47717 => x"00", -- $0ba65
          47718 => x"00", -- $0ba66
          47719 => x"00", -- $0ba67
          47720 => x"00", -- $0ba68
          47721 => x"00", -- $0ba69
          47722 => x"00", -- $0ba6a
          47723 => x"00", -- $0ba6b
          47724 => x"00", -- $0ba6c
          47725 => x"00", -- $0ba6d
          47726 => x"00", -- $0ba6e
          47727 => x"00", -- $0ba6f
          47728 => x"00", -- $0ba70
          47729 => x"00", -- $0ba71
          47730 => x"00", -- $0ba72
          47731 => x"00", -- $0ba73
          47732 => x"00", -- $0ba74
          47733 => x"00", -- $0ba75
          47734 => x"00", -- $0ba76
          47735 => x"00", -- $0ba77
          47736 => x"00", -- $0ba78
          47737 => x"00", -- $0ba79
          47738 => x"00", -- $0ba7a
          47739 => x"00", -- $0ba7b
          47740 => x"00", -- $0ba7c
          47741 => x"00", -- $0ba7d
          47742 => x"00", -- $0ba7e
          47743 => x"00", -- $0ba7f
          47744 => x"00", -- $0ba80
          47745 => x"00", -- $0ba81
          47746 => x"00", -- $0ba82
          47747 => x"00", -- $0ba83
          47748 => x"00", -- $0ba84
          47749 => x"00", -- $0ba85
          47750 => x"00", -- $0ba86
          47751 => x"00", -- $0ba87
          47752 => x"00", -- $0ba88
          47753 => x"00", -- $0ba89
          47754 => x"00", -- $0ba8a
          47755 => x"00", -- $0ba8b
          47756 => x"00", -- $0ba8c
          47757 => x"00", -- $0ba8d
          47758 => x"00", -- $0ba8e
          47759 => x"00", -- $0ba8f
          47760 => x"00", -- $0ba90
          47761 => x"00", -- $0ba91
          47762 => x"00", -- $0ba92
          47763 => x"00", -- $0ba93
          47764 => x"00", -- $0ba94
          47765 => x"00", -- $0ba95
          47766 => x"00", -- $0ba96
          47767 => x"00", -- $0ba97
          47768 => x"00", -- $0ba98
          47769 => x"00", -- $0ba99
          47770 => x"00", -- $0ba9a
          47771 => x"00", -- $0ba9b
          47772 => x"00", -- $0ba9c
          47773 => x"00", -- $0ba9d
          47774 => x"00", -- $0ba9e
          47775 => x"00", -- $0ba9f
          47776 => x"00", -- $0baa0
          47777 => x"00", -- $0baa1
          47778 => x"00", -- $0baa2
          47779 => x"00", -- $0baa3
          47780 => x"00", -- $0baa4
          47781 => x"00", -- $0baa5
          47782 => x"00", -- $0baa6
          47783 => x"00", -- $0baa7
          47784 => x"00", -- $0baa8
          47785 => x"00", -- $0baa9
          47786 => x"00", -- $0baaa
          47787 => x"00", -- $0baab
          47788 => x"00", -- $0baac
          47789 => x"00", -- $0baad
          47790 => x"00", -- $0baae
          47791 => x"00", -- $0baaf
          47792 => x"00", -- $0bab0
          47793 => x"00", -- $0bab1
          47794 => x"00", -- $0bab2
          47795 => x"00", -- $0bab3
          47796 => x"00", -- $0bab4
          47797 => x"00", -- $0bab5
          47798 => x"00", -- $0bab6
          47799 => x"00", -- $0bab7
          47800 => x"00", -- $0bab8
          47801 => x"00", -- $0bab9
          47802 => x"00", -- $0baba
          47803 => x"00", -- $0babb
          47804 => x"00", -- $0babc
          47805 => x"00", -- $0babd
          47806 => x"00", -- $0babe
          47807 => x"00", -- $0babf
          47808 => x"00", -- $0bac0
          47809 => x"00", -- $0bac1
          47810 => x"00", -- $0bac2
          47811 => x"00", -- $0bac3
          47812 => x"00", -- $0bac4
          47813 => x"00", -- $0bac5
          47814 => x"00", -- $0bac6
          47815 => x"00", -- $0bac7
          47816 => x"00", -- $0bac8
          47817 => x"00", -- $0bac9
          47818 => x"00", -- $0baca
          47819 => x"00", -- $0bacb
          47820 => x"00", -- $0bacc
          47821 => x"00", -- $0bacd
          47822 => x"00", -- $0bace
          47823 => x"00", -- $0bacf
          47824 => x"00", -- $0bad0
          47825 => x"00", -- $0bad1
          47826 => x"00", -- $0bad2
          47827 => x"00", -- $0bad3
          47828 => x"00", -- $0bad4
          47829 => x"00", -- $0bad5
          47830 => x"00", -- $0bad6
          47831 => x"00", -- $0bad7
          47832 => x"00", -- $0bad8
          47833 => x"00", -- $0bad9
          47834 => x"00", -- $0bada
          47835 => x"00", -- $0badb
          47836 => x"00", -- $0badc
          47837 => x"00", -- $0badd
          47838 => x"00", -- $0bade
          47839 => x"00", -- $0badf
          47840 => x"00", -- $0bae0
          47841 => x"00", -- $0bae1
          47842 => x"00", -- $0bae2
          47843 => x"00", -- $0bae3
          47844 => x"00", -- $0bae4
          47845 => x"00", -- $0bae5
          47846 => x"00", -- $0bae6
          47847 => x"00", -- $0bae7
          47848 => x"00", -- $0bae8
          47849 => x"00", -- $0bae9
          47850 => x"00", -- $0baea
          47851 => x"00", -- $0baeb
          47852 => x"00", -- $0baec
          47853 => x"00", -- $0baed
          47854 => x"00", -- $0baee
          47855 => x"00", -- $0baef
          47856 => x"00", -- $0baf0
          47857 => x"00", -- $0baf1
          47858 => x"00", -- $0baf2
          47859 => x"00", -- $0baf3
          47860 => x"00", -- $0baf4
          47861 => x"00", -- $0baf5
          47862 => x"00", -- $0baf6
          47863 => x"00", -- $0baf7
          47864 => x"00", -- $0baf8
          47865 => x"00", -- $0baf9
          47866 => x"00", -- $0bafa
          47867 => x"00", -- $0bafb
          47868 => x"00", -- $0bafc
          47869 => x"00", -- $0bafd
          47870 => x"00", -- $0bafe
          47871 => x"00", -- $0baff
          47872 => x"00", -- $0bb00
          47873 => x"00", -- $0bb01
          47874 => x"00", -- $0bb02
          47875 => x"00", -- $0bb03
          47876 => x"00", -- $0bb04
          47877 => x"00", -- $0bb05
          47878 => x"00", -- $0bb06
          47879 => x"00", -- $0bb07
          47880 => x"00", -- $0bb08
          47881 => x"00", -- $0bb09
          47882 => x"00", -- $0bb0a
          47883 => x"00", -- $0bb0b
          47884 => x"00", -- $0bb0c
          47885 => x"00", -- $0bb0d
          47886 => x"00", -- $0bb0e
          47887 => x"00", -- $0bb0f
          47888 => x"00", -- $0bb10
          47889 => x"00", -- $0bb11
          47890 => x"00", -- $0bb12
          47891 => x"00", -- $0bb13
          47892 => x"00", -- $0bb14
          47893 => x"00", -- $0bb15
          47894 => x"00", -- $0bb16
          47895 => x"00", -- $0bb17
          47896 => x"00", -- $0bb18
          47897 => x"00", -- $0bb19
          47898 => x"00", -- $0bb1a
          47899 => x"00", -- $0bb1b
          47900 => x"00", -- $0bb1c
          47901 => x"00", -- $0bb1d
          47902 => x"00", -- $0bb1e
          47903 => x"00", -- $0bb1f
          47904 => x"00", -- $0bb20
          47905 => x"00", -- $0bb21
          47906 => x"00", -- $0bb22
          47907 => x"00", -- $0bb23
          47908 => x"00", -- $0bb24
          47909 => x"00", -- $0bb25
          47910 => x"00", -- $0bb26
          47911 => x"00", -- $0bb27
          47912 => x"00", -- $0bb28
          47913 => x"00", -- $0bb29
          47914 => x"00", -- $0bb2a
          47915 => x"00", -- $0bb2b
          47916 => x"00", -- $0bb2c
          47917 => x"00", -- $0bb2d
          47918 => x"00", -- $0bb2e
          47919 => x"00", -- $0bb2f
          47920 => x"00", -- $0bb30
          47921 => x"00", -- $0bb31
          47922 => x"00", -- $0bb32
          47923 => x"00", -- $0bb33
          47924 => x"00", -- $0bb34
          47925 => x"00", -- $0bb35
          47926 => x"00", -- $0bb36
          47927 => x"00", -- $0bb37
          47928 => x"00", -- $0bb38
          47929 => x"00", -- $0bb39
          47930 => x"00", -- $0bb3a
          47931 => x"00", -- $0bb3b
          47932 => x"00", -- $0bb3c
          47933 => x"00", -- $0bb3d
          47934 => x"00", -- $0bb3e
          47935 => x"00", -- $0bb3f
          47936 => x"00", -- $0bb40
          47937 => x"00", -- $0bb41
          47938 => x"00", -- $0bb42
          47939 => x"00", -- $0bb43
          47940 => x"00", -- $0bb44
          47941 => x"00", -- $0bb45
          47942 => x"00", -- $0bb46
          47943 => x"00", -- $0bb47
          47944 => x"00", -- $0bb48
          47945 => x"00", -- $0bb49
          47946 => x"00", -- $0bb4a
          47947 => x"00", -- $0bb4b
          47948 => x"00", -- $0bb4c
          47949 => x"00", -- $0bb4d
          47950 => x"00", -- $0bb4e
          47951 => x"00", -- $0bb4f
          47952 => x"00", -- $0bb50
          47953 => x"00", -- $0bb51
          47954 => x"00", -- $0bb52
          47955 => x"00", -- $0bb53
          47956 => x"00", -- $0bb54
          47957 => x"00", -- $0bb55
          47958 => x"00", -- $0bb56
          47959 => x"00", -- $0bb57
          47960 => x"00", -- $0bb58
          47961 => x"00", -- $0bb59
          47962 => x"00", -- $0bb5a
          47963 => x"00", -- $0bb5b
          47964 => x"00", -- $0bb5c
          47965 => x"00", -- $0bb5d
          47966 => x"00", -- $0bb5e
          47967 => x"00", -- $0bb5f
          47968 => x"00", -- $0bb60
          47969 => x"00", -- $0bb61
          47970 => x"00", -- $0bb62
          47971 => x"00", -- $0bb63
          47972 => x"00", -- $0bb64
          47973 => x"00", -- $0bb65
          47974 => x"00", -- $0bb66
          47975 => x"00", -- $0bb67
          47976 => x"00", -- $0bb68
          47977 => x"00", -- $0bb69
          47978 => x"00", -- $0bb6a
          47979 => x"00", -- $0bb6b
          47980 => x"00", -- $0bb6c
          47981 => x"00", -- $0bb6d
          47982 => x"00", -- $0bb6e
          47983 => x"00", -- $0bb6f
          47984 => x"00", -- $0bb70
          47985 => x"00", -- $0bb71
          47986 => x"00", -- $0bb72
          47987 => x"00", -- $0bb73
          47988 => x"00", -- $0bb74
          47989 => x"00", -- $0bb75
          47990 => x"00", -- $0bb76
          47991 => x"00", -- $0bb77
          47992 => x"00", -- $0bb78
          47993 => x"00", -- $0bb79
          47994 => x"00", -- $0bb7a
          47995 => x"00", -- $0bb7b
          47996 => x"00", -- $0bb7c
          47997 => x"00", -- $0bb7d
          47998 => x"00", -- $0bb7e
          47999 => x"00", -- $0bb7f
          48000 => x"00", -- $0bb80
          48001 => x"00", -- $0bb81
          48002 => x"00", -- $0bb82
          48003 => x"00", -- $0bb83
          48004 => x"00", -- $0bb84
          48005 => x"00", -- $0bb85
          48006 => x"00", -- $0bb86
          48007 => x"00", -- $0bb87
          48008 => x"00", -- $0bb88
          48009 => x"00", -- $0bb89
          48010 => x"00", -- $0bb8a
          48011 => x"00", -- $0bb8b
          48012 => x"00", -- $0bb8c
          48013 => x"00", -- $0bb8d
          48014 => x"00", -- $0bb8e
          48015 => x"00", -- $0bb8f
          48016 => x"00", -- $0bb90
          48017 => x"00", -- $0bb91
          48018 => x"00", -- $0bb92
          48019 => x"00", -- $0bb93
          48020 => x"00", -- $0bb94
          48021 => x"00", -- $0bb95
          48022 => x"00", -- $0bb96
          48023 => x"00", -- $0bb97
          48024 => x"00", -- $0bb98
          48025 => x"00", -- $0bb99
          48026 => x"00", -- $0bb9a
          48027 => x"00", -- $0bb9b
          48028 => x"00", -- $0bb9c
          48029 => x"00", -- $0bb9d
          48030 => x"00", -- $0bb9e
          48031 => x"00", -- $0bb9f
          48032 => x"00", -- $0bba0
          48033 => x"00", -- $0bba1
          48034 => x"00", -- $0bba2
          48035 => x"00", -- $0bba3
          48036 => x"00", -- $0bba4
          48037 => x"00", -- $0bba5
          48038 => x"00", -- $0bba6
          48039 => x"00", -- $0bba7
          48040 => x"00", -- $0bba8
          48041 => x"00", -- $0bba9
          48042 => x"00", -- $0bbaa
          48043 => x"00", -- $0bbab
          48044 => x"00", -- $0bbac
          48045 => x"00", -- $0bbad
          48046 => x"00", -- $0bbae
          48047 => x"00", -- $0bbaf
          48048 => x"00", -- $0bbb0
          48049 => x"00", -- $0bbb1
          48050 => x"00", -- $0bbb2
          48051 => x"00", -- $0bbb3
          48052 => x"00", -- $0bbb4
          48053 => x"00", -- $0bbb5
          48054 => x"00", -- $0bbb6
          48055 => x"00", -- $0bbb7
          48056 => x"00", -- $0bbb8
          48057 => x"00", -- $0bbb9
          48058 => x"00", -- $0bbba
          48059 => x"00", -- $0bbbb
          48060 => x"00", -- $0bbbc
          48061 => x"00", -- $0bbbd
          48062 => x"00", -- $0bbbe
          48063 => x"00", -- $0bbbf
          48064 => x"00", -- $0bbc0
          48065 => x"00", -- $0bbc1
          48066 => x"00", -- $0bbc2
          48067 => x"00", -- $0bbc3
          48068 => x"00", -- $0bbc4
          48069 => x"00", -- $0bbc5
          48070 => x"00", -- $0bbc6
          48071 => x"00", -- $0bbc7
          48072 => x"00", -- $0bbc8
          48073 => x"00", -- $0bbc9
          48074 => x"00", -- $0bbca
          48075 => x"00", -- $0bbcb
          48076 => x"00", -- $0bbcc
          48077 => x"00", -- $0bbcd
          48078 => x"00", -- $0bbce
          48079 => x"00", -- $0bbcf
          48080 => x"00", -- $0bbd0
          48081 => x"00", -- $0bbd1
          48082 => x"00", -- $0bbd2
          48083 => x"00", -- $0bbd3
          48084 => x"00", -- $0bbd4
          48085 => x"00", -- $0bbd5
          48086 => x"00", -- $0bbd6
          48087 => x"00", -- $0bbd7
          48088 => x"00", -- $0bbd8
          48089 => x"00", -- $0bbd9
          48090 => x"00", -- $0bbda
          48091 => x"00", -- $0bbdb
          48092 => x"00", -- $0bbdc
          48093 => x"00", -- $0bbdd
          48094 => x"00", -- $0bbde
          48095 => x"00", -- $0bbdf
          48096 => x"00", -- $0bbe0
          48097 => x"00", -- $0bbe1
          48098 => x"00", -- $0bbe2
          48099 => x"00", -- $0bbe3
          48100 => x"00", -- $0bbe4
          48101 => x"00", -- $0bbe5
          48102 => x"00", -- $0bbe6
          48103 => x"00", -- $0bbe7
          48104 => x"00", -- $0bbe8
          48105 => x"00", -- $0bbe9
          48106 => x"00", -- $0bbea
          48107 => x"00", -- $0bbeb
          48108 => x"00", -- $0bbec
          48109 => x"00", -- $0bbed
          48110 => x"00", -- $0bbee
          48111 => x"00", -- $0bbef
          48112 => x"00", -- $0bbf0
          48113 => x"00", -- $0bbf1
          48114 => x"00", -- $0bbf2
          48115 => x"00", -- $0bbf3
          48116 => x"00", -- $0bbf4
          48117 => x"00", -- $0bbf5
          48118 => x"00", -- $0bbf6
          48119 => x"00", -- $0bbf7
          48120 => x"00", -- $0bbf8
          48121 => x"00", -- $0bbf9
          48122 => x"00", -- $0bbfa
          48123 => x"00", -- $0bbfb
          48124 => x"00", -- $0bbfc
          48125 => x"00", -- $0bbfd
          48126 => x"00", -- $0bbfe
          48127 => x"00", -- $0bbff
          48128 => x"00", -- $0bc00
          48129 => x"00", -- $0bc01
          48130 => x"00", -- $0bc02
          48131 => x"00", -- $0bc03
          48132 => x"00", -- $0bc04
          48133 => x"00", -- $0bc05
          48134 => x"00", -- $0bc06
          48135 => x"00", -- $0bc07
          48136 => x"00", -- $0bc08
          48137 => x"00", -- $0bc09
          48138 => x"00", -- $0bc0a
          48139 => x"00", -- $0bc0b
          48140 => x"00", -- $0bc0c
          48141 => x"00", -- $0bc0d
          48142 => x"00", -- $0bc0e
          48143 => x"00", -- $0bc0f
          48144 => x"00", -- $0bc10
          48145 => x"00", -- $0bc11
          48146 => x"00", -- $0bc12
          48147 => x"00", -- $0bc13
          48148 => x"00", -- $0bc14
          48149 => x"00", -- $0bc15
          48150 => x"00", -- $0bc16
          48151 => x"00", -- $0bc17
          48152 => x"00", -- $0bc18
          48153 => x"00", -- $0bc19
          48154 => x"00", -- $0bc1a
          48155 => x"00", -- $0bc1b
          48156 => x"00", -- $0bc1c
          48157 => x"00", -- $0bc1d
          48158 => x"00", -- $0bc1e
          48159 => x"00", -- $0bc1f
          48160 => x"00", -- $0bc20
          48161 => x"00", -- $0bc21
          48162 => x"00", -- $0bc22
          48163 => x"00", -- $0bc23
          48164 => x"00", -- $0bc24
          48165 => x"00", -- $0bc25
          48166 => x"00", -- $0bc26
          48167 => x"00", -- $0bc27
          48168 => x"00", -- $0bc28
          48169 => x"00", -- $0bc29
          48170 => x"00", -- $0bc2a
          48171 => x"00", -- $0bc2b
          48172 => x"00", -- $0bc2c
          48173 => x"00", -- $0bc2d
          48174 => x"00", -- $0bc2e
          48175 => x"00", -- $0bc2f
          48176 => x"00", -- $0bc30
          48177 => x"00", -- $0bc31
          48178 => x"00", -- $0bc32
          48179 => x"00", -- $0bc33
          48180 => x"00", -- $0bc34
          48181 => x"00", -- $0bc35
          48182 => x"00", -- $0bc36
          48183 => x"00", -- $0bc37
          48184 => x"00", -- $0bc38
          48185 => x"00", -- $0bc39
          48186 => x"00", -- $0bc3a
          48187 => x"00", -- $0bc3b
          48188 => x"00", -- $0bc3c
          48189 => x"00", -- $0bc3d
          48190 => x"00", -- $0bc3e
          48191 => x"00", -- $0bc3f
          48192 => x"00", -- $0bc40
          48193 => x"00", -- $0bc41
          48194 => x"00", -- $0bc42
          48195 => x"00", -- $0bc43
          48196 => x"00", -- $0bc44
          48197 => x"00", -- $0bc45
          48198 => x"00", -- $0bc46
          48199 => x"00", -- $0bc47
          48200 => x"00", -- $0bc48
          48201 => x"00", -- $0bc49
          48202 => x"00", -- $0bc4a
          48203 => x"00", -- $0bc4b
          48204 => x"00", -- $0bc4c
          48205 => x"00", -- $0bc4d
          48206 => x"00", -- $0bc4e
          48207 => x"00", -- $0bc4f
          48208 => x"00", -- $0bc50
          48209 => x"00", -- $0bc51
          48210 => x"00", -- $0bc52
          48211 => x"00", -- $0bc53
          48212 => x"00", -- $0bc54
          48213 => x"00", -- $0bc55
          48214 => x"00", -- $0bc56
          48215 => x"00", -- $0bc57
          48216 => x"00", -- $0bc58
          48217 => x"00", -- $0bc59
          48218 => x"00", -- $0bc5a
          48219 => x"00", -- $0bc5b
          48220 => x"00", -- $0bc5c
          48221 => x"00", -- $0bc5d
          48222 => x"00", -- $0bc5e
          48223 => x"00", -- $0bc5f
          48224 => x"00", -- $0bc60
          48225 => x"00", -- $0bc61
          48226 => x"00", -- $0bc62
          48227 => x"00", -- $0bc63
          48228 => x"00", -- $0bc64
          48229 => x"00", -- $0bc65
          48230 => x"00", -- $0bc66
          48231 => x"00", -- $0bc67
          48232 => x"00", -- $0bc68
          48233 => x"00", -- $0bc69
          48234 => x"00", -- $0bc6a
          48235 => x"00", -- $0bc6b
          48236 => x"00", -- $0bc6c
          48237 => x"00", -- $0bc6d
          48238 => x"00", -- $0bc6e
          48239 => x"00", -- $0bc6f
          48240 => x"00", -- $0bc70
          48241 => x"00", -- $0bc71
          48242 => x"00", -- $0bc72
          48243 => x"00", -- $0bc73
          48244 => x"00", -- $0bc74
          48245 => x"00", -- $0bc75
          48246 => x"00", -- $0bc76
          48247 => x"00", -- $0bc77
          48248 => x"00", -- $0bc78
          48249 => x"00", -- $0bc79
          48250 => x"00", -- $0bc7a
          48251 => x"00", -- $0bc7b
          48252 => x"00", -- $0bc7c
          48253 => x"00", -- $0bc7d
          48254 => x"00", -- $0bc7e
          48255 => x"00", -- $0bc7f
          48256 => x"00", -- $0bc80
          48257 => x"00", -- $0bc81
          48258 => x"00", -- $0bc82
          48259 => x"00", -- $0bc83
          48260 => x"00", -- $0bc84
          48261 => x"00", -- $0bc85
          48262 => x"00", -- $0bc86
          48263 => x"00", -- $0bc87
          48264 => x"00", -- $0bc88
          48265 => x"00", -- $0bc89
          48266 => x"00", -- $0bc8a
          48267 => x"00", -- $0bc8b
          48268 => x"00", -- $0bc8c
          48269 => x"00", -- $0bc8d
          48270 => x"00", -- $0bc8e
          48271 => x"00", -- $0bc8f
          48272 => x"00", -- $0bc90
          48273 => x"00", -- $0bc91
          48274 => x"00", -- $0bc92
          48275 => x"00", -- $0bc93
          48276 => x"00", -- $0bc94
          48277 => x"00", -- $0bc95
          48278 => x"00", -- $0bc96
          48279 => x"00", -- $0bc97
          48280 => x"00", -- $0bc98
          48281 => x"00", -- $0bc99
          48282 => x"00", -- $0bc9a
          48283 => x"00", -- $0bc9b
          48284 => x"00", -- $0bc9c
          48285 => x"00", -- $0bc9d
          48286 => x"00", -- $0bc9e
          48287 => x"00", -- $0bc9f
          48288 => x"00", -- $0bca0
          48289 => x"00", -- $0bca1
          48290 => x"00", -- $0bca2
          48291 => x"00", -- $0bca3
          48292 => x"00", -- $0bca4
          48293 => x"00", -- $0bca5
          48294 => x"00", -- $0bca6
          48295 => x"00", -- $0bca7
          48296 => x"00", -- $0bca8
          48297 => x"00", -- $0bca9
          48298 => x"00", -- $0bcaa
          48299 => x"00", -- $0bcab
          48300 => x"00", -- $0bcac
          48301 => x"00", -- $0bcad
          48302 => x"00", -- $0bcae
          48303 => x"00", -- $0bcaf
          48304 => x"00", -- $0bcb0
          48305 => x"00", -- $0bcb1
          48306 => x"00", -- $0bcb2
          48307 => x"00", -- $0bcb3
          48308 => x"00", -- $0bcb4
          48309 => x"00", -- $0bcb5
          48310 => x"00", -- $0bcb6
          48311 => x"00", -- $0bcb7
          48312 => x"00", -- $0bcb8
          48313 => x"00", -- $0bcb9
          48314 => x"00", -- $0bcba
          48315 => x"00", -- $0bcbb
          48316 => x"00", -- $0bcbc
          48317 => x"00", -- $0bcbd
          48318 => x"00", -- $0bcbe
          48319 => x"00", -- $0bcbf
          48320 => x"00", -- $0bcc0
          48321 => x"00", -- $0bcc1
          48322 => x"00", -- $0bcc2
          48323 => x"00", -- $0bcc3
          48324 => x"00", -- $0bcc4
          48325 => x"00", -- $0bcc5
          48326 => x"00", -- $0bcc6
          48327 => x"00", -- $0bcc7
          48328 => x"00", -- $0bcc8
          48329 => x"00", -- $0bcc9
          48330 => x"00", -- $0bcca
          48331 => x"00", -- $0bccb
          48332 => x"00", -- $0bccc
          48333 => x"00", -- $0bccd
          48334 => x"00", -- $0bcce
          48335 => x"00", -- $0bccf
          48336 => x"00", -- $0bcd0
          48337 => x"00", -- $0bcd1
          48338 => x"00", -- $0bcd2
          48339 => x"00", -- $0bcd3
          48340 => x"00", -- $0bcd4
          48341 => x"00", -- $0bcd5
          48342 => x"00", -- $0bcd6
          48343 => x"00", -- $0bcd7
          48344 => x"00", -- $0bcd8
          48345 => x"00", -- $0bcd9
          48346 => x"00", -- $0bcda
          48347 => x"00", -- $0bcdb
          48348 => x"00", -- $0bcdc
          48349 => x"00", -- $0bcdd
          48350 => x"00", -- $0bcde
          48351 => x"00", -- $0bcdf
          48352 => x"00", -- $0bce0
          48353 => x"00", -- $0bce1
          48354 => x"00", -- $0bce2
          48355 => x"00", -- $0bce3
          48356 => x"00", -- $0bce4
          48357 => x"00", -- $0bce5
          48358 => x"00", -- $0bce6
          48359 => x"00", -- $0bce7
          48360 => x"00", -- $0bce8
          48361 => x"00", -- $0bce9
          48362 => x"00", -- $0bcea
          48363 => x"00", -- $0bceb
          48364 => x"00", -- $0bcec
          48365 => x"00", -- $0bced
          48366 => x"00", -- $0bcee
          48367 => x"00", -- $0bcef
          48368 => x"00", -- $0bcf0
          48369 => x"00", -- $0bcf1
          48370 => x"00", -- $0bcf2
          48371 => x"00", -- $0bcf3
          48372 => x"00", -- $0bcf4
          48373 => x"00", -- $0bcf5
          48374 => x"00", -- $0bcf6
          48375 => x"00", -- $0bcf7
          48376 => x"00", -- $0bcf8
          48377 => x"00", -- $0bcf9
          48378 => x"00", -- $0bcfa
          48379 => x"00", -- $0bcfb
          48380 => x"00", -- $0bcfc
          48381 => x"00", -- $0bcfd
          48382 => x"00", -- $0bcfe
          48383 => x"00", -- $0bcff
          48384 => x"00", -- $0bd00
          48385 => x"00", -- $0bd01
          48386 => x"00", -- $0bd02
          48387 => x"00", -- $0bd03
          48388 => x"00", -- $0bd04
          48389 => x"00", -- $0bd05
          48390 => x"00", -- $0bd06
          48391 => x"00", -- $0bd07
          48392 => x"00", -- $0bd08
          48393 => x"00", -- $0bd09
          48394 => x"00", -- $0bd0a
          48395 => x"00", -- $0bd0b
          48396 => x"00", -- $0bd0c
          48397 => x"00", -- $0bd0d
          48398 => x"00", -- $0bd0e
          48399 => x"00", -- $0bd0f
          48400 => x"00", -- $0bd10
          48401 => x"00", -- $0bd11
          48402 => x"00", -- $0bd12
          48403 => x"00", -- $0bd13
          48404 => x"00", -- $0bd14
          48405 => x"00", -- $0bd15
          48406 => x"00", -- $0bd16
          48407 => x"00", -- $0bd17
          48408 => x"00", -- $0bd18
          48409 => x"00", -- $0bd19
          48410 => x"00", -- $0bd1a
          48411 => x"00", -- $0bd1b
          48412 => x"00", -- $0bd1c
          48413 => x"00", -- $0bd1d
          48414 => x"00", -- $0bd1e
          48415 => x"00", -- $0bd1f
          48416 => x"00", -- $0bd20
          48417 => x"00", -- $0bd21
          48418 => x"00", -- $0bd22
          48419 => x"00", -- $0bd23
          48420 => x"00", -- $0bd24
          48421 => x"00", -- $0bd25
          48422 => x"00", -- $0bd26
          48423 => x"00", -- $0bd27
          48424 => x"00", -- $0bd28
          48425 => x"00", -- $0bd29
          48426 => x"00", -- $0bd2a
          48427 => x"00", -- $0bd2b
          48428 => x"00", -- $0bd2c
          48429 => x"00", -- $0bd2d
          48430 => x"00", -- $0bd2e
          48431 => x"00", -- $0bd2f
          48432 => x"00", -- $0bd30
          48433 => x"00", -- $0bd31
          48434 => x"00", -- $0bd32
          48435 => x"00", -- $0bd33
          48436 => x"00", -- $0bd34
          48437 => x"00", -- $0bd35
          48438 => x"00", -- $0bd36
          48439 => x"00", -- $0bd37
          48440 => x"00", -- $0bd38
          48441 => x"00", -- $0bd39
          48442 => x"00", -- $0bd3a
          48443 => x"00", -- $0bd3b
          48444 => x"00", -- $0bd3c
          48445 => x"00", -- $0bd3d
          48446 => x"00", -- $0bd3e
          48447 => x"00", -- $0bd3f
          48448 => x"00", -- $0bd40
          48449 => x"00", -- $0bd41
          48450 => x"00", -- $0bd42
          48451 => x"00", -- $0bd43
          48452 => x"00", -- $0bd44
          48453 => x"00", -- $0bd45
          48454 => x"00", -- $0bd46
          48455 => x"00", -- $0bd47
          48456 => x"00", -- $0bd48
          48457 => x"00", -- $0bd49
          48458 => x"00", -- $0bd4a
          48459 => x"00", -- $0bd4b
          48460 => x"00", -- $0bd4c
          48461 => x"00", -- $0bd4d
          48462 => x"00", -- $0bd4e
          48463 => x"00", -- $0bd4f
          48464 => x"00", -- $0bd50
          48465 => x"00", -- $0bd51
          48466 => x"00", -- $0bd52
          48467 => x"00", -- $0bd53
          48468 => x"00", -- $0bd54
          48469 => x"00", -- $0bd55
          48470 => x"00", -- $0bd56
          48471 => x"00", -- $0bd57
          48472 => x"00", -- $0bd58
          48473 => x"00", -- $0bd59
          48474 => x"00", -- $0bd5a
          48475 => x"00", -- $0bd5b
          48476 => x"00", -- $0bd5c
          48477 => x"00", -- $0bd5d
          48478 => x"00", -- $0bd5e
          48479 => x"00", -- $0bd5f
          48480 => x"00", -- $0bd60
          48481 => x"00", -- $0bd61
          48482 => x"00", -- $0bd62
          48483 => x"00", -- $0bd63
          48484 => x"00", -- $0bd64
          48485 => x"00", -- $0bd65
          48486 => x"00", -- $0bd66
          48487 => x"00", -- $0bd67
          48488 => x"00", -- $0bd68
          48489 => x"00", -- $0bd69
          48490 => x"00", -- $0bd6a
          48491 => x"00", -- $0bd6b
          48492 => x"00", -- $0bd6c
          48493 => x"00", -- $0bd6d
          48494 => x"00", -- $0bd6e
          48495 => x"00", -- $0bd6f
          48496 => x"00", -- $0bd70
          48497 => x"00", -- $0bd71
          48498 => x"00", -- $0bd72
          48499 => x"00", -- $0bd73
          48500 => x"00", -- $0bd74
          48501 => x"00", -- $0bd75
          48502 => x"00", -- $0bd76
          48503 => x"00", -- $0bd77
          48504 => x"00", -- $0bd78
          48505 => x"00", -- $0bd79
          48506 => x"00", -- $0bd7a
          48507 => x"00", -- $0bd7b
          48508 => x"00", -- $0bd7c
          48509 => x"00", -- $0bd7d
          48510 => x"00", -- $0bd7e
          48511 => x"00", -- $0bd7f
          48512 => x"00", -- $0bd80
          48513 => x"00", -- $0bd81
          48514 => x"00", -- $0bd82
          48515 => x"00", -- $0bd83
          48516 => x"00", -- $0bd84
          48517 => x"00", -- $0bd85
          48518 => x"00", -- $0bd86
          48519 => x"00", -- $0bd87
          48520 => x"00", -- $0bd88
          48521 => x"00", -- $0bd89
          48522 => x"00", -- $0bd8a
          48523 => x"00", -- $0bd8b
          48524 => x"00", -- $0bd8c
          48525 => x"00", -- $0bd8d
          48526 => x"00", -- $0bd8e
          48527 => x"00", -- $0bd8f
          48528 => x"00", -- $0bd90
          48529 => x"00", -- $0bd91
          48530 => x"00", -- $0bd92
          48531 => x"00", -- $0bd93
          48532 => x"00", -- $0bd94
          48533 => x"00", -- $0bd95
          48534 => x"00", -- $0bd96
          48535 => x"00", -- $0bd97
          48536 => x"00", -- $0bd98
          48537 => x"00", -- $0bd99
          48538 => x"00", -- $0bd9a
          48539 => x"00", -- $0bd9b
          48540 => x"00", -- $0bd9c
          48541 => x"00", -- $0bd9d
          48542 => x"00", -- $0bd9e
          48543 => x"00", -- $0bd9f
          48544 => x"00", -- $0bda0
          48545 => x"00", -- $0bda1
          48546 => x"00", -- $0bda2
          48547 => x"00", -- $0bda3
          48548 => x"00", -- $0bda4
          48549 => x"00", -- $0bda5
          48550 => x"00", -- $0bda6
          48551 => x"00", -- $0bda7
          48552 => x"00", -- $0bda8
          48553 => x"00", -- $0bda9
          48554 => x"00", -- $0bdaa
          48555 => x"00", -- $0bdab
          48556 => x"00", -- $0bdac
          48557 => x"00", -- $0bdad
          48558 => x"00", -- $0bdae
          48559 => x"00", -- $0bdaf
          48560 => x"00", -- $0bdb0
          48561 => x"00", -- $0bdb1
          48562 => x"00", -- $0bdb2
          48563 => x"00", -- $0bdb3
          48564 => x"00", -- $0bdb4
          48565 => x"00", -- $0bdb5
          48566 => x"00", -- $0bdb6
          48567 => x"00", -- $0bdb7
          48568 => x"00", -- $0bdb8
          48569 => x"00", -- $0bdb9
          48570 => x"00", -- $0bdba
          48571 => x"00", -- $0bdbb
          48572 => x"00", -- $0bdbc
          48573 => x"00", -- $0bdbd
          48574 => x"00", -- $0bdbe
          48575 => x"00", -- $0bdbf
          48576 => x"00", -- $0bdc0
          48577 => x"00", -- $0bdc1
          48578 => x"00", -- $0bdc2
          48579 => x"00", -- $0bdc3
          48580 => x"00", -- $0bdc4
          48581 => x"00", -- $0bdc5
          48582 => x"00", -- $0bdc6
          48583 => x"00", -- $0bdc7
          48584 => x"00", -- $0bdc8
          48585 => x"00", -- $0bdc9
          48586 => x"00", -- $0bdca
          48587 => x"00", -- $0bdcb
          48588 => x"00", -- $0bdcc
          48589 => x"00", -- $0bdcd
          48590 => x"00", -- $0bdce
          48591 => x"00", -- $0bdcf
          48592 => x"00", -- $0bdd0
          48593 => x"00", -- $0bdd1
          48594 => x"00", -- $0bdd2
          48595 => x"00", -- $0bdd3
          48596 => x"00", -- $0bdd4
          48597 => x"00", -- $0bdd5
          48598 => x"00", -- $0bdd6
          48599 => x"00", -- $0bdd7
          48600 => x"00", -- $0bdd8
          48601 => x"00", -- $0bdd9
          48602 => x"00", -- $0bdda
          48603 => x"00", -- $0bddb
          48604 => x"00", -- $0bddc
          48605 => x"00", -- $0bddd
          48606 => x"00", -- $0bdde
          48607 => x"00", -- $0bddf
          48608 => x"00", -- $0bde0
          48609 => x"00", -- $0bde1
          48610 => x"00", -- $0bde2
          48611 => x"00", -- $0bde3
          48612 => x"00", -- $0bde4
          48613 => x"00", -- $0bde5
          48614 => x"00", -- $0bde6
          48615 => x"00", -- $0bde7
          48616 => x"00", -- $0bde8
          48617 => x"00", -- $0bde9
          48618 => x"00", -- $0bdea
          48619 => x"00", -- $0bdeb
          48620 => x"00", -- $0bdec
          48621 => x"00", -- $0bded
          48622 => x"00", -- $0bdee
          48623 => x"00", -- $0bdef
          48624 => x"00", -- $0bdf0
          48625 => x"00", -- $0bdf1
          48626 => x"00", -- $0bdf2
          48627 => x"00", -- $0bdf3
          48628 => x"00", -- $0bdf4
          48629 => x"00", -- $0bdf5
          48630 => x"00", -- $0bdf6
          48631 => x"00", -- $0bdf7
          48632 => x"00", -- $0bdf8
          48633 => x"00", -- $0bdf9
          48634 => x"00", -- $0bdfa
          48635 => x"00", -- $0bdfb
          48636 => x"00", -- $0bdfc
          48637 => x"00", -- $0bdfd
          48638 => x"00", -- $0bdfe
          48639 => x"00", -- $0bdff
          48640 => x"00", -- $0be00
          48641 => x"00", -- $0be01
          48642 => x"00", -- $0be02
          48643 => x"00", -- $0be03
          48644 => x"00", -- $0be04
          48645 => x"00", -- $0be05
          48646 => x"00", -- $0be06
          48647 => x"00", -- $0be07
          48648 => x"00", -- $0be08
          48649 => x"00", -- $0be09
          48650 => x"00", -- $0be0a
          48651 => x"00", -- $0be0b
          48652 => x"00", -- $0be0c
          48653 => x"00", -- $0be0d
          48654 => x"00", -- $0be0e
          48655 => x"00", -- $0be0f
          48656 => x"00", -- $0be10
          48657 => x"00", -- $0be11
          48658 => x"00", -- $0be12
          48659 => x"00", -- $0be13
          48660 => x"00", -- $0be14
          48661 => x"00", -- $0be15
          48662 => x"00", -- $0be16
          48663 => x"00", -- $0be17
          48664 => x"00", -- $0be18
          48665 => x"00", -- $0be19
          48666 => x"00", -- $0be1a
          48667 => x"00", -- $0be1b
          48668 => x"00", -- $0be1c
          48669 => x"00", -- $0be1d
          48670 => x"00", -- $0be1e
          48671 => x"00", -- $0be1f
          48672 => x"00", -- $0be20
          48673 => x"00", -- $0be21
          48674 => x"00", -- $0be22
          48675 => x"00", -- $0be23
          48676 => x"00", -- $0be24
          48677 => x"00", -- $0be25
          48678 => x"00", -- $0be26
          48679 => x"00", -- $0be27
          48680 => x"00", -- $0be28
          48681 => x"00", -- $0be29
          48682 => x"00", -- $0be2a
          48683 => x"00", -- $0be2b
          48684 => x"00", -- $0be2c
          48685 => x"00", -- $0be2d
          48686 => x"00", -- $0be2e
          48687 => x"00", -- $0be2f
          48688 => x"00", -- $0be30
          48689 => x"00", -- $0be31
          48690 => x"00", -- $0be32
          48691 => x"00", -- $0be33
          48692 => x"00", -- $0be34
          48693 => x"00", -- $0be35
          48694 => x"00", -- $0be36
          48695 => x"00", -- $0be37
          48696 => x"00", -- $0be38
          48697 => x"00", -- $0be39
          48698 => x"00", -- $0be3a
          48699 => x"00", -- $0be3b
          48700 => x"00", -- $0be3c
          48701 => x"00", -- $0be3d
          48702 => x"00", -- $0be3e
          48703 => x"00", -- $0be3f
          48704 => x"00", -- $0be40
          48705 => x"00", -- $0be41
          48706 => x"00", -- $0be42
          48707 => x"00", -- $0be43
          48708 => x"00", -- $0be44
          48709 => x"00", -- $0be45
          48710 => x"00", -- $0be46
          48711 => x"00", -- $0be47
          48712 => x"00", -- $0be48
          48713 => x"00", -- $0be49
          48714 => x"00", -- $0be4a
          48715 => x"00", -- $0be4b
          48716 => x"00", -- $0be4c
          48717 => x"00", -- $0be4d
          48718 => x"00", -- $0be4e
          48719 => x"00", -- $0be4f
          48720 => x"00", -- $0be50
          48721 => x"00", -- $0be51
          48722 => x"00", -- $0be52
          48723 => x"00", -- $0be53
          48724 => x"00", -- $0be54
          48725 => x"00", -- $0be55
          48726 => x"00", -- $0be56
          48727 => x"00", -- $0be57
          48728 => x"00", -- $0be58
          48729 => x"00", -- $0be59
          48730 => x"00", -- $0be5a
          48731 => x"00", -- $0be5b
          48732 => x"00", -- $0be5c
          48733 => x"00", -- $0be5d
          48734 => x"00", -- $0be5e
          48735 => x"00", -- $0be5f
          48736 => x"00", -- $0be60
          48737 => x"00", -- $0be61
          48738 => x"00", -- $0be62
          48739 => x"00", -- $0be63
          48740 => x"00", -- $0be64
          48741 => x"00", -- $0be65
          48742 => x"00", -- $0be66
          48743 => x"00", -- $0be67
          48744 => x"00", -- $0be68
          48745 => x"00", -- $0be69
          48746 => x"00", -- $0be6a
          48747 => x"00", -- $0be6b
          48748 => x"00", -- $0be6c
          48749 => x"00", -- $0be6d
          48750 => x"00", -- $0be6e
          48751 => x"00", -- $0be6f
          48752 => x"00", -- $0be70
          48753 => x"00", -- $0be71
          48754 => x"00", -- $0be72
          48755 => x"00", -- $0be73
          48756 => x"00", -- $0be74
          48757 => x"00", -- $0be75
          48758 => x"00", -- $0be76
          48759 => x"00", -- $0be77
          48760 => x"00", -- $0be78
          48761 => x"00", -- $0be79
          48762 => x"00", -- $0be7a
          48763 => x"00", -- $0be7b
          48764 => x"00", -- $0be7c
          48765 => x"00", -- $0be7d
          48766 => x"00", -- $0be7e
          48767 => x"00", -- $0be7f
          48768 => x"00", -- $0be80
          48769 => x"00", -- $0be81
          48770 => x"00", -- $0be82
          48771 => x"00", -- $0be83
          48772 => x"00", -- $0be84
          48773 => x"00", -- $0be85
          48774 => x"00", -- $0be86
          48775 => x"00", -- $0be87
          48776 => x"00", -- $0be88
          48777 => x"00", -- $0be89
          48778 => x"00", -- $0be8a
          48779 => x"00", -- $0be8b
          48780 => x"00", -- $0be8c
          48781 => x"00", -- $0be8d
          48782 => x"00", -- $0be8e
          48783 => x"00", -- $0be8f
          48784 => x"00", -- $0be90
          48785 => x"00", -- $0be91
          48786 => x"00", -- $0be92
          48787 => x"00", -- $0be93
          48788 => x"00", -- $0be94
          48789 => x"00", -- $0be95
          48790 => x"00", -- $0be96
          48791 => x"00", -- $0be97
          48792 => x"00", -- $0be98
          48793 => x"00", -- $0be99
          48794 => x"00", -- $0be9a
          48795 => x"00", -- $0be9b
          48796 => x"00", -- $0be9c
          48797 => x"00", -- $0be9d
          48798 => x"00", -- $0be9e
          48799 => x"00", -- $0be9f
          48800 => x"00", -- $0bea0
          48801 => x"00", -- $0bea1
          48802 => x"00", -- $0bea2
          48803 => x"00", -- $0bea3
          48804 => x"00", -- $0bea4
          48805 => x"00", -- $0bea5
          48806 => x"00", -- $0bea6
          48807 => x"00", -- $0bea7
          48808 => x"00", -- $0bea8
          48809 => x"00", -- $0bea9
          48810 => x"00", -- $0beaa
          48811 => x"00", -- $0beab
          48812 => x"00", -- $0beac
          48813 => x"00", -- $0bead
          48814 => x"00", -- $0beae
          48815 => x"00", -- $0beaf
          48816 => x"00", -- $0beb0
          48817 => x"00", -- $0beb1
          48818 => x"00", -- $0beb2
          48819 => x"00", -- $0beb3
          48820 => x"00", -- $0beb4
          48821 => x"00", -- $0beb5
          48822 => x"00", -- $0beb6
          48823 => x"00", -- $0beb7
          48824 => x"00", -- $0beb8
          48825 => x"00", -- $0beb9
          48826 => x"00", -- $0beba
          48827 => x"00", -- $0bebb
          48828 => x"00", -- $0bebc
          48829 => x"00", -- $0bebd
          48830 => x"00", -- $0bebe
          48831 => x"00", -- $0bebf
          48832 => x"00", -- $0bec0
          48833 => x"00", -- $0bec1
          48834 => x"00", -- $0bec2
          48835 => x"00", -- $0bec3
          48836 => x"00", -- $0bec4
          48837 => x"00", -- $0bec5
          48838 => x"00", -- $0bec6
          48839 => x"00", -- $0bec7
          48840 => x"00", -- $0bec8
          48841 => x"00", -- $0bec9
          48842 => x"00", -- $0beca
          48843 => x"00", -- $0becb
          48844 => x"00", -- $0becc
          48845 => x"00", -- $0becd
          48846 => x"00", -- $0bece
          48847 => x"00", -- $0becf
          48848 => x"00", -- $0bed0
          48849 => x"00", -- $0bed1
          48850 => x"00", -- $0bed2
          48851 => x"00", -- $0bed3
          48852 => x"00", -- $0bed4
          48853 => x"00", -- $0bed5
          48854 => x"00", -- $0bed6
          48855 => x"00", -- $0bed7
          48856 => x"00", -- $0bed8
          48857 => x"00", -- $0bed9
          48858 => x"00", -- $0beda
          48859 => x"00", -- $0bedb
          48860 => x"00", -- $0bedc
          48861 => x"00", -- $0bedd
          48862 => x"00", -- $0bede
          48863 => x"00", -- $0bedf
          48864 => x"00", -- $0bee0
          48865 => x"00", -- $0bee1
          48866 => x"00", -- $0bee2
          48867 => x"00", -- $0bee3
          48868 => x"00", -- $0bee4
          48869 => x"00", -- $0bee5
          48870 => x"00", -- $0bee6
          48871 => x"00", -- $0bee7
          48872 => x"00", -- $0bee8
          48873 => x"00", -- $0bee9
          48874 => x"00", -- $0beea
          48875 => x"00", -- $0beeb
          48876 => x"00", -- $0beec
          48877 => x"00", -- $0beed
          48878 => x"00", -- $0beee
          48879 => x"00", -- $0beef
          48880 => x"00", -- $0bef0
          48881 => x"00", -- $0bef1
          48882 => x"00", -- $0bef2
          48883 => x"00", -- $0bef3
          48884 => x"00", -- $0bef4
          48885 => x"00", -- $0bef5
          48886 => x"00", -- $0bef6
          48887 => x"00", -- $0bef7
          48888 => x"00", -- $0bef8
          48889 => x"00", -- $0bef9
          48890 => x"00", -- $0befa
          48891 => x"00", -- $0befb
          48892 => x"00", -- $0befc
          48893 => x"00", -- $0befd
          48894 => x"00", -- $0befe
          48895 => x"00", -- $0beff
          48896 => x"00", -- $0bf00
          48897 => x"00", -- $0bf01
          48898 => x"00", -- $0bf02
          48899 => x"00", -- $0bf03
          48900 => x"00", -- $0bf04
          48901 => x"00", -- $0bf05
          48902 => x"00", -- $0bf06
          48903 => x"00", -- $0bf07
          48904 => x"00", -- $0bf08
          48905 => x"00", -- $0bf09
          48906 => x"00", -- $0bf0a
          48907 => x"00", -- $0bf0b
          48908 => x"00", -- $0bf0c
          48909 => x"00", -- $0bf0d
          48910 => x"00", -- $0bf0e
          48911 => x"00", -- $0bf0f
          48912 => x"00", -- $0bf10
          48913 => x"00", -- $0bf11
          48914 => x"00", -- $0bf12
          48915 => x"00", -- $0bf13
          48916 => x"00", -- $0bf14
          48917 => x"00", -- $0bf15
          48918 => x"00", -- $0bf16
          48919 => x"00", -- $0bf17
          48920 => x"00", -- $0bf18
          48921 => x"00", -- $0bf19
          48922 => x"00", -- $0bf1a
          48923 => x"00", -- $0bf1b
          48924 => x"00", -- $0bf1c
          48925 => x"00", -- $0bf1d
          48926 => x"00", -- $0bf1e
          48927 => x"00", -- $0bf1f
          48928 => x"00", -- $0bf20
          48929 => x"00", -- $0bf21
          48930 => x"00", -- $0bf22
          48931 => x"00", -- $0bf23
          48932 => x"00", -- $0bf24
          48933 => x"00", -- $0bf25
          48934 => x"00", -- $0bf26
          48935 => x"00", -- $0bf27
          48936 => x"00", -- $0bf28
          48937 => x"00", -- $0bf29
          48938 => x"00", -- $0bf2a
          48939 => x"00", -- $0bf2b
          48940 => x"00", -- $0bf2c
          48941 => x"00", -- $0bf2d
          48942 => x"00", -- $0bf2e
          48943 => x"00", -- $0bf2f
          48944 => x"00", -- $0bf30
          48945 => x"00", -- $0bf31
          48946 => x"00", -- $0bf32
          48947 => x"00", -- $0bf33
          48948 => x"00", -- $0bf34
          48949 => x"00", -- $0bf35
          48950 => x"00", -- $0bf36
          48951 => x"00", -- $0bf37
          48952 => x"00", -- $0bf38
          48953 => x"00", -- $0bf39
          48954 => x"00", -- $0bf3a
          48955 => x"00", -- $0bf3b
          48956 => x"00", -- $0bf3c
          48957 => x"00", -- $0bf3d
          48958 => x"00", -- $0bf3e
          48959 => x"00", -- $0bf3f
          48960 => x"00", -- $0bf40
          48961 => x"00", -- $0bf41
          48962 => x"00", -- $0bf42
          48963 => x"00", -- $0bf43
          48964 => x"00", -- $0bf44
          48965 => x"00", -- $0bf45
          48966 => x"00", -- $0bf46
          48967 => x"00", -- $0bf47
          48968 => x"00", -- $0bf48
          48969 => x"00", -- $0bf49
          48970 => x"00", -- $0bf4a
          48971 => x"00", -- $0bf4b
          48972 => x"00", -- $0bf4c
          48973 => x"00", -- $0bf4d
          48974 => x"00", -- $0bf4e
          48975 => x"00", -- $0bf4f
          48976 => x"00", -- $0bf50
          48977 => x"00", -- $0bf51
          48978 => x"00", -- $0bf52
          48979 => x"00", -- $0bf53
          48980 => x"00", -- $0bf54
          48981 => x"00", -- $0bf55
          48982 => x"00", -- $0bf56
          48983 => x"00", -- $0bf57
          48984 => x"00", -- $0bf58
          48985 => x"00", -- $0bf59
          48986 => x"00", -- $0bf5a
          48987 => x"00", -- $0bf5b
          48988 => x"00", -- $0bf5c
          48989 => x"00", -- $0bf5d
          48990 => x"00", -- $0bf5e
          48991 => x"00", -- $0bf5f
          48992 => x"00", -- $0bf60
          48993 => x"00", -- $0bf61
          48994 => x"00", -- $0bf62
          48995 => x"00", -- $0bf63
          48996 => x"00", -- $0bf64
          48997 => x"00", -- $0bf65
          48998 => x"00", -- $0bf66
          48999 => x"00", -- $0bf67
          49000 => x"00", -- $0bf68
          49001 => x"00", -- $0bf69
          49002 => x"00", -- $0bf6a
          49003 => x"00", -- $0bf6b
          49004 => x"00", -- $0bf6c
          49005 => x"00", -- $0bf6d
          49006 => x"00", -- $0bf6e
          49007 => x"00", -- $0bf6f
          49008 => x"00", -- $0bf70
          49009 => x"00", -- $0bf71
          49010 => x"00", -- $0bf72
          49011 => x"00", -- $0bf73
          49012 => x"00", -- $0bf74
          49013 => x"00", -- $0bf75
          49014 => x"00", -- $0bf76
          49015 => x"00", -- $0bf77
          49016 => x"00", -- $0bf78
          49017 => x"00", -- $0bf79
          49018 => x"00", -- $0bf7a
          49019 => x"00", -- $0bf7b
          49020 => x"00", -- $0bf7c
          49021 => x"00", -- $0bf7d
          49022 => x"00", -- $0bf7e
          49023 => x"00", -- $0bf7f
          49024 => x"00", -- $0bf80
          49025 => x"00", -- $0bf81
          49026 => x"00", -- $0bf82
          49027 => x"00", -- $0bf83
          49028 => x"00", -- $0bf84
          49029 => x"00", -- $0bf85
          49030 => x"00", -- $0bf86
          49031 => x"00", -- $0bf87
          49032 => x"00", -- $0bf88
          49033 => x"00", -- $0bf89
          49034 => x"00", -- $0bf8a
          49035 => x"00", -- $0bf8b
          49036 => x"00", -- $0bf8c
          49037 => x"00", -- $0bf8d
          49038 => x"00", -- $0bf8e
          49039 => x"00", -- $0bf8f
          49040 => x"00", -- $0bf90
          49041 => x"00", -- $0bf91
          49042 => x"00", -- $0bf92
          49043 => x"00", -- $0bf93
          49044 => x"00", -- $0bf94
          49045 => x"00", -- $0bf95
          49046 => x"00", -- $0bf96
          49047 => x"00", -- $0bf97
          49048 => x"00", -- $0bf98
          49049 => x"00", -- $0bf99
          49050 => x"00", -- $0bf9a
          49051 => x"00", -- $0bf9b
          49052 => x"00", -- $0bf9c
          49053 => x"00", -- $0bf9d
          49054 => x"00", -- $0bf9e
          49055 => x"00", -- $0bf9f
          49056 => x"00", -- $0bfa0
          49057 => x"00", -- $0bfa1
          49058 => x"00", -- $0bfa2
          49059 => x"00", -- $0bfa3
          49060 => x"00", -- $0bfa4
          49061 => x"00", -- $0bfa5
          49062 => x"00", -- $0bfa6
          49063 => x"00", -- $0bfa7
          49064 => x"00", -- $0bfa8
          49065 => x"00", -- $0bfa9
          49066 => x"00", -- $0bfaa
          49067 => x"00", -- $0bfab
          49068 => x"00", -- $0bfac
          49069 => x"00", -- $0bfad
          49070 => x"00", -- $0bfae
          49071 => x"00", -- $0bfaf
          49072 => x"00", -- $0bfb0
          49073 => x"00", -- $0bfb1
          49074 => x"00", -- $0bfb2
          49075 => x"00", -- $0bfb3
          49076 => x"00", -- $0bfb4
          49077 => x"00", -- $0bfb5
          49078 => x"00", -- $0bfb6
          49079 => x"00", -- $0bfb7
          49080 => x"00", -- $0bfb8
          49081 => x"00", -- $0bfb9
          49082 => x"00", -- $0bfba
          49083 => x"00", -- $0bfbb
          49084 => x"00", -- $0bfbc
          49085 => x"00", -- $0bfbd
          49086 => x"00", -- $0bfbe
          49087 => x"00", -- $0bfbf
          49088 => x"00", -- $0bfc0
          49089 => x"00", -- $0bfc1
          49090 => x"00", -- $0bfc2
          49091 => x"00", -- $0bfc3
          49092 => x"00", -- $0bfc4
          49093 => x"00", -- $0bfc5
          49094 => x"00", -- $0bfc6
          49095 => x"00", -- $0bfc7
          49096 => x"00", -- $0bfc8
          49097 => x"00", -- $0bfc9
          49098 => x"00", -- $0bfca
          49099 => x"00", -- $0bfcb
          49100 => x"00", -- $0bfcc
          49101 => x"00", -- $0bfcd
          49102 => x"00", -- $0bfce
          49103 => x"00", -- $0bfcf
          49104 => x"00", -- $0bfd0
          49105 => x"00", -- $0bfd1
          49106 => x"00", -- $0bfd2
          49107 => x"00", -- $0bfd3
          49108 => x"00", -- $0bfd4
          49109 => x"00", -- $0bfd5
          49110 => x"00", -- $0bfd6
          49111 => x"00", -- $0bfd7
          49112 => x"00", -- $0bfd8
          49113 => x"00", -- $0bfd9
          49114 => x"00", -- $0bfda
          49115 => x"00", -- $0bfdb
          49116 => x"00", -- $0bfdc
          49117 => x"00", -- $0bfdd
          49118 => x"00", -- $0bfde
          49119 => x"00", -- $0bfdf
          49120 => x"00", -- $0bfe0
          49121 => x"00", -- $0bfe1
          49122 => x"00", -- $0bfe2
          49123 => x"00", -- $0bfe3
          49124 => x"00", -- $0bfe4
          49125 => x"00", -- $0bfe5
          49126 => x"00", -- $0bfe6
          49127 => x"00", -- $0bfe7
          49128 => x"00", -- $0bfe8
          49129 => x"00", -- $0bfe9
          49130 => x"00", -- $0bfea
          49131 => x"00", -- $0bfeb
          49132 => x"00", -- $0bfec
          49133 => x"00", -- $0bfed
          49134 => x"00", -- $0bfee
          49135 => x"00", -- $0bfef
          49136 => x"00", -- $0bff0
          49137 => x"00", -- $0bff1
          49138 => x"00", -- $0bff2
          49139 => x"00", -- $0bff3
          49140 => x"00", -- $0bff4
          49141 => x"00", -- $0bff5
          49142 => x"00", -- $0bff6
          49143 => x"00", -- $0bff7
          49144 => x"00", -- $0bff8
          49145 => x"00", -- $0bff9
          49146 => x"00", -- $0bffa
          49147 => x"00", -- $0bffb
          49148 => x"00", -- $0bffc
          49149 => x"00", -- $0bffd
          49150 => x"00", -- $0bffe
          49151 => x"00", -- $0bfff
          49152 => x"00", -- $0c000
          49153 => x"00", -- $0c001
          49154 => x"00", -- $0c002
          49155 => x"00", -- $0c003
          49156 => x"00", -- $0c004
          49157 => x"00", -- $0c005
          49158 => x"00", -- $0c006
          49159 => x"00", -- $0c007
          49160 => x"00", -- $0c008
          49161 => x"00", -- $0c009
          49162 => x"00", -- $0c00a
          49163 => x"00", -- $0c00b
          49164 => x"00", -- $0c00c
          49165 => x"00", -- $0c00d
          49166 => x"00", -- $0c00e
          49167 => x"00", -- $0c00f
          49168 => x"00", -- $0c010
          49169 => x"00", -- $0c011
          49170 => x"00", -- $0c012
          49171 => x"00", -- $0c013
          49172 => x"00", -- $0c014
          49173 => x"00", -- $0c015
          49174 => x"00", -- $0c016
          49175 => x"00", -- $0c017
          49176 => x"00", -- $0c018
          49177 => x"00", -- $0c019
          49178 => x"00", -- $0c01a
          49179 => x"00", -- $0c01b
          49180 => x"00", -- $0c01c
          49181 => x"00", -- $0c01d
          49182 => x"00", -- $0c01e
          49183 => x"00", -- $0c01f
          49184 => x"00", -- $0c020
          49185 => x"00", -- $0c021
          49186 => x"00", -- $0c022
          49187 => x"00", -- $0c023
          49188 => x"00", -- $0c024
          49189 => x"00", -- $0c025
          49190 => x"00", -- $0c026
          49191 => x"00", -- $0c027
          49192 => x"00", -- $0c028
          49193 => x"00", -- $0c029
          49194 => x"00", -- $0c02a
          49195 => x"00", -- $0c02b
          49196 => x"00", -- $0c02c
          49197 => x"00", -- $0c02d
          49198 => x"00", -- $0c02e
          49199 => x"00", -- $0c02f
          49200 => x"00", -- $0c030
          49201 => x"00", -- $0c031
          49202 => x"00", -- $0c032
          49203 => x"00", -- $0c033
          49204 => x"00", -- $0c034
          49205 => x"00", -- $0c035
          49206 => x"00", -- $0c036
          49207 => x"00", -- $0c037
          49208 => x"00", -- $0c038
          49209 => x"00", -- $0c039
          49210 => x"00", -- $0c03a
          49211 => x"00", -- $0c03b
          49212 => x"00", -- $0c03c
          49213 => x"00", -- $0c03d
          49214 => x"00", -- $0c03e
          49215 => x"00", -- $0c03f
          49216 => x"00", -- $0c040
          49217 => x"00", -- $0c041
          49218 => x"00", -- $0c042
          49219 => x"00", -- $0c043
          49220 => x"00", -- $0c044
          49221 => x"00", -- $0c045
          49222 => x"00", -- $0c046
          49223 => x"00", -- $0c047
          49224 => x"00", -- $0c048
          49225 => x"00", -- $0c049
          49226 => x"00", -- $0c04a
          49227 => x"00", -- $0c04b
          49228 => x"00", -- $0c04c
          49229 => x"00", -- $0c04d
          49230 => x"00", -- $0c04e
          49231 => x"00", -- $0c04f
          49232 => x"00", -- $0c050
          49233 => x"00", -- $0c051
          49234 => x"00", -- $0c052
          49235 => x"00", -- $0c053
          49236 => x"00", -- $0c054
          49237 => x"00", -- $0c055
          49238 => x"00", -- $0c056
          49239 => x"00", -- $0c057
          49240 => x"00", -- $0c058
          49241 => x"00", -- $0c059
          49242 => x"00", -- $0c05a
          49243 => x"00", -- $0c05b
          49244 => x"00", -- $0c05c
          49245 => x"00", -- $0c05d
          49246 => x"00", -- $0c05e
          49247 => x"00", -- $0c05f
          49248 => x"00", -- $0c060
          49249 => x"00", -- $0c061
          49250 => x"00", -- $0c062
          49251 => x"00", -- $0c063
          49252 => x"00", -- $0c064
          49253 => x"00", -- $0c065
          49254 => x"00", -- $0c066
          49255 => x"00", -- $0c067
          49256 => x"00", -- $0c068
          49257 => x"00", -- $0c069
          49258 => x"00", -- $0c06a
          49259 => x"00", -- $0c06b
          49260 => x"00", -- $0c06c
          49261 => x"00", -- $0c06d
          49262 => x"00", -- $0c06e
          49263 => x"00", -- $0c06f
          49264 => x"00", -- $0c070
          49265 => x"00", -- $0c071
          49266 => x"00", -- $0c072
          49267 => x"00", -- $0c073
          49268 => x"00", -- $0c074
          49269 => x"00", -- $0c075
          49270 => x"00", -- $0c076
          49271 => x"00", -- $0c077
          49272 => x"00", -- $0c078
          49273 => x"00", -- $0c079
          49274 => x"00", -- $0c07a
          49275 => x"00", -- $0c07b
          49276 => x"00", -- $0c07c
          49277 => x"00", -- $0c07d
          49278 => x"00", -- $0c07e
          49279 => x"00", -- $0c07f
          49280 => x"00", -- $0c080
          49281 => x"00", -- $0c081
          49282 => x"00", -- $0c082
          49283 => x"00", -- $0c083
          49284 => x"00", -- $0c084
          49285 => x"00", -- $0c085
          49286 => x"00", -- $0c086
          49287 => x"00", -- $0c087
          49288 => x"00", -- $0c088
          49289 => x"00", -- $0c089
          49290 => x"00", -- $0c08a
          49291 => x"00", -- $0c08b
          49292 => x"00", -- $0c08c
          49293 => x"00", -- $0c08d
          49294 => x"00", -- $0c08e
          49295 => x"00", -- $0c08f
          49296 => x"00", -- $0c090
          49297 => x"00", -- $0c091
          49298 => x"00", -- $0c092
          49299 => x"00", -- $0c093
          49300 => x"00", -- $0c094
          49301 => x"00", -- $0c095
          49302 => x"00", -- $0c096
          49303 => x"00", -- $0c097
          49304 => x"00", -- $0c098
          49305 => x"00", -- $0c099
          49306 => x"00", -- $0c09a
          49307 => x"00", -- $0c09b
          49308 => x"00", -- $0c09c
          49309 => x"00", -- $0c09d
          49310 => x"00", -- $0c09e
          49311 => x"00", -- $0c09f
          49312 => x"00", -- $0c0a0
          49313 => x"00", -- $0c0a1
          49314 => x"00", -- $0c0a2
          49315 => x"00", -- $0c0a3
          49316 => x"00", -- $0c0a4
          49317 => x"00", -- $0c0a5
          49318 => x"00", -- $0c0a6
          49319 => x"00", -- $0c0a7
          49320 => x"00", -- $0c0a8
          49321 => x"00", -- $0c0a9
          49322 => x"00", -- $0c0aa
          49323 => x"00", -- $0c0ab
          49324 => x"00", -- $0c0ac
          49325 => x"00", -- $0c0ad
          49326 => x"00", -- $0c0ae
          49327 => x"00", -- $0c0af
          49328 => x"00", -- $0c0b0
          49329 => x"00", -- $0c0b1
          49330 => x"00", -- $0c0b2
          49331 => x"00", -- $0c0b3
          49332 => x"00", -- $0c0b4
          49333 => x"00", -- $0c0b5
          49334 => x"00", -- $0c0b6
          49335 => x"00", -- $0c0b7
          49336 => x"00", -- $0c0b8
          49337 => x"00", -- $0c0b9
          49338 => x"00", -- $0c0ba
          49339 => x"00", -- $0c0bb
          49340 => x"00", -- $0c0bc
          49341 => x"00", -- $0c0bd
          49342 => x"00", -- $0c0be
          49343 => x"00", -- $0c0bf
          49344 => x"00", -- $0c0c0
          49345 => x"00", -- $0c0c1
          49346 => x"00", -- $0c0c2
          49347 => x"00", -- $0c0c3
          49348 => x"00", -- $0c0c4
          49349 => x"00", -- $0c0c5
          49350 => x"00", -- $0c0c6
          49351 => x"00", -- $0c0c7
          49352 => x"00", -- $0c0c8
          49353 => x"00", -- $0c0c9
          49354 => x"00", -- $0c0ca
          49355 => x"00", -- $0c0cb
          49356 => x"00", -- $0c0cc
          49357 => x"00", -- $0c0cd
          49358 => x"00", -- $0c0ce
          49359 => x"00", -- $0c0cf
          49360 => x"00", -- $0c0d0
          49361 => x"00", -- $0c0d1
          49362 => x"00", -- $0c0d2
          49363 => x"00", -- $0c0d3
          49364 => x"00", -- $0c0d4
          49365 => x"00", -- $0c0d5
          49366 => x"00", -- $0c0d6
          49367 => x"00", -- $0c0d7
          49368 => x"00", -- $0c0d8
          49369 => x"00", -- $0c0d9
          49370 => x"00", -- $0c0da
          49371 => x"00", -- $0c0db
          49372 => x"00", -- $0c0dc
          49373 => x"00", -- $0c0dd
          49374 => x"00", -- $0c0de
          49375 => x"00", -- $0c0df
          49376 => x"00", -- $0c0e0
          49377 => x"00", -- $0c0e1
          49378 => x"00", -- $0c0e2
          49379 => x"00", -- $0c0e3
          49380 => x"00", -- $0c0e4
          49381 => x"00", -- $0c0e5
          49382 => x"00", -- $0c0e6
          49383 => x"00", -- $0c0e7
          49384 => x"00", -- $0c0e8
          49385 => x"00", -- $0c0e9
          49386 => x"00", -- $0c0ea
          49387 => x"00", -- $0c0eb
          49388 => x"00", -- $0c0ec
          49389 => x"00", -- $0c0ed
          49390 => x"00", -- $0c0ee
          49391 => x"00", -- $0c0ef
          49392 => x"00", -- $0c0f0
          49393 => x"00", -- $0c0f1
          49394 => x"00", -- $0c0f2
          49395 => x"00", -- $0c0f3
          49396 => x"00", -- $0c0f4
          49397 => x"00", -- $0c0f5
          49398 => x"00", -- $0c0f6
          49399 => x"00", -- $0c0f7
          49400 => x"00", -- $0c0f8
          49401 => x"00", -- $0c0f9
          49402 => x"00", -- $0c0fa
          49403 => x"00", -- $0c0fb
          49404 => x"00", -- $0c0fc
          49405 => x"00", -- $0c0fd
          49406 => x"00", -- $0c0fe
          49407 => x"00", -- $0c0ff
          49408 => x"00", -- $0c100
          49409 => x"00", -- $0c101
          49410 => x"00", -- $0c102
          49411 => x"00", -- $0c103
          49412 => x"00", -- $0c104
          49413 => x"00", -- $0c105
          49414 => x"00", -- $0c106
          49415 => x"00", -- $0c107
          49416 => x"00", -- $0c108
          49417 => x"00", -- $0c109
          49418 => x"00", -- $0c10a
          49419 => x"00", -- $0c10b
          49420 => x"00", -- $0c10c
          49421 => x"00", -- $0c10d
          49422 => x"00", -- $0c10e
          49423 => x"00", -- $0c10f
          49424 => x"00", -- $0c110
          49425 => x"00", -- $0c111
          49426 => x"00", -- $0c112
          49427 => x"00", -- $0c113
          49428 => x"00", -- $0c114
          49429 => x"00", -- $0c115
          49430 => x"00", -- $0c116
          49431 => x"00", -- $0c117
          49432 => x"00", -- $0c118
          49433 => x"00", -- $0c119
          49434 => x"00", -- $0c11a
          49435 => x"00", -- $0c11b
          49436 => x"00", -- $0c11c
          49437 => x"00", -- $0c11d
          49438 => x"00", -- $0c11e
          49439 => x"00", -- $0c11f
          49440 => x"00", -- $0c120
          49441 => x"00", -- $0c121
          49442 => x"00", -- $0c122
          49443 => x"00", -- $0c123
          49444 => x"00", -- $0c124
          49445 => x"00", -- $0c125
          49446 => x"00", -- $0c126
          49447 => x"00", -- $0c127
          49448 => x"00", -- $0c128
          49449 => x"00", -- $0c129
          49450 => x"00", -- $0c12a
          49451 => x"00", -- $0c12b
          49452 => x"00", -- $0c12c
          49453 => x"00", -- $0c12d
          49454 => x"00", -- $0c12e
          49455 => x"00", -- $0c12f
          49456 => x"00", -- $0c130
          49457 => x"00", -- $0c131
          49458 => x"00", -- $0c132
          49459 => x"00", -- $0c133
          49460 => x"00", -- $0c134
          49461 => x"00", -- $0c135
          49462 => x"00", -- $0c136
          49463 => x"00", -- $0c137
          49464 => x"00", -- $0c138
          49465 => x"00", -- $0c139
          49466 => x"00", -- $0c13a
          49467 => x"00", -- $0c13b
          49468 => x"00", -- $0c13c
          49469 => x"00", -- $0c13d
          49470 => x"00", -- $0c13e
          49471 => x"00", -- $0c13f
          49472 => x"00", -- $0c140
          49473 => x"00", -- $0c141
          49474 => x"00", -- $0c142
          49475 => x"00", -- $0c143
          49476 => x"00", -- $0c144
          49477 => x"00", -- $0c145
          49478 => x"00", -- $0c146
          49479 => x"00", -- $0c147
          49480 => x"00", -- $0c148
          49481 => x"00", -- $0c149
          49482 => x"00", -- $0c14a
          49483 => x"00", -- $0c14b
          49484 => x"00", -- $0c14c
          49485 => x"00", -- $0c14d
          49486 => x"00", -- $0c14e
          49487 => x"00", -- $0c14f
          49488 => x"00", -- $0c150
          49489 => x"00", -- $0c151
          49490 => x"00", -- $0c152
          49491 => x"00", -- $0c153
          49492 => x"00", -- $0c154
          49493 => x"00", -- $0c155
          49494 => x"00", -- $0c156
          49495 => x"00", -- $0c157
          49496 => x"00", -- $0c158
          49497 => x"00", -- $0c159
          49498 => x"00", -- $0c15a
          49499 => x"00", -- $0c15b
          49500 => x"00", -- $0c15c
          49501 => x"00", -- $0c15d
          49502 => x"00", -- $0c15e
          49503 => x"00", -- $0c15f
          49504 => x"00", -- $0c160
          49505 => x"00", -- $0c161
          49506 => x"00", -- $0c162
          49507 => x"00", -- $0c163
          49508 => x"00", -- $0c164
          49509 => x"00", -- $0c165
          49510 => x"00", -- $0c166
          49511 => x"00", -- $0c167
          49512 => x"00", -- $0c168
          49513 => x"00", -- $0c169
          49514 => x"00", -- $0c16a
          49515 => x"00", -- $0c16b
          49516 => x"00", -- $0c16c
          49517 => x"00", -- $0c16d
          49518 => x"00", -- $0c16e
          49519 => x"00", -- $0c16f
          49520 => x"00", -- $0c170
          49521 => x"00", -- $0c171
          49522 => x"00", -- $0c172
          49523 => x"00", -- $0c173
          49524 => x"00", -- $0c174
          49525 => x"00", -- $0c175
          49526 => x"00", -- $0c176
          49527 => x"00", -- $0c177
          49528 => x"00", -- $0c178
          49529 => x"00", -- $0c179
          49530 => x"00", -- $0c17a
          49531 => x"00", -- $0c17b
          49532 => x"00", -- $0c17c
          49533 => x"00", -- $0c17d
          49534 => x"00", -- $0c17e
          49535 => x"00", -- $0c17f
          49536 => x"00", -- $0c180
          49537 => x"00", -- $0c181
          49538 => x"00", -- $0c182
          49539 => x"00", -- $0c183
          49540 => x"00", -- $0c184
          49541 => x"00", -- $0c185
          49542 => x"00", -- $0c186
          49543 => x"00", -- $0c187
          49544 => x"00", -- $0c188
          49545 => x"00", -- $0c189
          49546 => x"00", -- $0c18a
          49547 => x"00", -- $0c18b
          49548 => x"00", -- $0c18c
          49549 => x"00", -- $0c18d
          49550 => x"00", -- $0c18e
          49551 => x"00", -- $0c18f
          49552 => x"00", -- $0c190
          49553 => x"00", -- $0c191
          49554 => x"00", -- $0c192
          49555 => x"00", -- $0c193
          49556 => x"00", -- $0c194
          49557 => x"00", -- $0c195
          49558 => x"00", -- $0c196
          49559 => x"00", -- $0c197
          49560 => x"00", -- $0c198
          49561 => x"00", -- $0c199
          49562 => x"00", -- $0c19a
          49563 => x"00", -- $0c19b
          49564 => x"00", -- $0c19c
          49565 => x"00", -- $0c19d
          49566 => x"00", -- $0c19e
          49567 => x"00", -- $0c19f
          49568 => x"00", -- $0c1a0
          49569 => x"00", -- $0c1a1
          49570 => x"00", -- $0c1a2
          49571 => x"00", -- $0c1a3
          49572 => x"00", -- $0c1a4
          49573 => x"00", -- $0c1a5
          49574 => x"00", -- $0c1a6
          49575 => x"00", -- $0c1a7
          49576 => x"00", -- $0c1a8
          49577 => x"00", -- $0c1a9
          49578 => x"00", -- $0c1aa
          49579 => x"00", -- $0c1ab
          49580 => x"00", -- $0c1ac
          49581 => x"00", -- $0c1ad
          49582 => x"00", -- $0c1ae
          49583 => x"00", -- $0c1af
          49584 => x"00", -- $0c1b0
          49585 => x"00", -- $0c1b1
          49586 => x"00", -- $0c1b2
          49587 => x"00", -- $0c1b3
          49588 => x"00", -- $0c1b4
          49589 => x"00", -- $0c1b5
          49590 => x"00", -- $0c1b6
          49591 => x"00", -- $0c1b7
          49592 => x"00", -- $0c1b8
          49593 => x"00", -- $0c1b9
          49594 => x"00", -- $0c1ba
          49595 => x"00", -- $0c1bb
          49596 => x"00", -- $0c1bc
          49597 => x"00", -- $0c1bd
          49598 => x"00", -- $0c1be
          49599 => x"00", -- $0c1bf
          49600 => x"00", -- $0c1c0
          49601 => x"00", -- $0c1c1
          49602 => x"00", -- $0c1c2
          49603 => x"00", -- $0c1c3
          49604 => x"00", -- $0c1c4
          49605 => x"00", -- $0c1c5
          49606 => x"00", -- $0c1c6
          49607 => x"00", -- $0c1c7
          49608 => x"00", -- $0c1c8
          49609 => x"00", -- $0c1c9
          49610 => x"00", -- $0c1ca
          49611 => x"00", -- $0c1cb
          49612 => x"00", -- $0c1cc
          49613 => x"00", -- $0c1cd
          49614 => x"00", -- $0c1ce
          49615 => x"00", -- $0c1cf
          49616 => x"00", -- $0c1d0
          49617 => x"00", -- $0c1d1
          49618 => x"00", -- $0c1d2
          49619 => x"00", -- $0c1d3
          49620 => x"00", -- $0c1d4
          49621 => x"00", -- $0c1d5
          49622 => x"00", -- $0c1d6
          49623 => x"00", -- $0c1d7
          49624 => x"00", -- $0c1d8
          49625 => x"00", -- $0c1d9
          49626 => x"00", -- $0c1da
          49627 => x"00", -- $0c1db
          49628 => x"00", -- $0c1dc
          49629 => x"00", -- $0c1dd
          49630 => x"00", -- $0c1de
          49631 => x"00", -- $0c1df
          49632 => x"00", -- $0c1e0
          49633 => x"00", -- $0c1e1
          49634 => x"00", -- $0c1e2
          49635 => x"00", -- $0c1e3
          49636 => x"00", -- $0c1e4
          49637 => x"00", -- $0c1e5
          49638 => x"00", -- $0c1e6
          49639 => x"00", -- $0c1e7
          49640 => x"00", -- $0c1e8
          49641 => x"00", -- $0c1e9
          49642 => x"00", -- $0c1ea
          49643 => x"00", -- $0c1eb
          49644 => x"00", -- $0c1ec
          49645 => x"00", -- $0c1ed
          49646 => x"00", -- $0c1ee
          49647 => x"00", -- $0c1ef
          49648 => x"00", -- $0c1f0
          49649 => x"00", -- $0c1f1
          49650 => x"00", -- $0c1f2
          49651 => x"00", -- $0c1f3
          49652 => x"00", -- $0c1f4
          49653 => x"00", -- $0c1f5
          49654 => x"00", -- $0c1f6
          49655 => x"00", -- $0c1f7
          49656 => x"00", -- $0c1f8
          49657 => x"00", -- $0c1f9
          49658 => x"00", -- $0c1fa
          49659 => x"00", -- $0c1fb
          49660 => x"00", -- $0c1fc
          49661 => x"00", -- $0c1fd
          49662 => x"00", -- $0c1fe
          49663 => x"00", -- $0c1ff
          49664 => x"00", -- $0c200
          49665 => x"00", -- $0c201
          49666 => x"00", -- $0c202
          49667 => x"00", -- $0c203
          49668 => x"00", -- $0c204
          49669 => x"00", -- $0c205
          49670 => x"00", -- $0c206
          49671 => x"00", -- $0c207
          49672 => x"00", -- $0c208
          49673 => x"00", -- $0c209
          49674 => x"00", -- $0c20a
          49675 => x"00", -- $0c20b
          49676 => x"00", -- $0c20c
          49677 => x"00", -- $0c20d
          49678 => x"00", -- $0c20e
          49679 => x"00", -- $0c20f
          49680 => x"00", -- $0c210
          49681 => x"00", -- $0c211
          49682 => x"00", -- $0c212
          49683 => x"00", -- $0c213
          49684 => x"00", -- $0c214
          49685 => x"00", -- $0c215
          49686 => x"00", -- $0c216
          49687 => x"00", -- $0c217
          49688 => x"00", -- $0c218
          49689 => x"00", -- $0c219
          49690 => x"00", -- $0c21a
          49691 => x"00", -- $0c21b
          49692 => x"00", -- $0c21c
          49693 => x"00", -- $0c21d
          49694 => x"00", -- $0c21e
          49695 => x"00", -- $0c21f
          49696 => x"00", -- $0c220
          49697 => x"00", -- $0c221
          49698 => x"00", -- $0c222
          49699 => x"00", -- $0c223
          49700 => x"00", -- $0c224
          49701 => x"00", -- $0c225
          49702 => x"00", -- $0c226
          49703 => x"00", -- $0c227
          49704 => x"00", -- $0c228
          49705 => x"00", -- $0c229
          49706 => x"00", -- $0c22a
          49707 => x"00", -- $0c22b
          49708 => x"00", -- $0c22c
          49709 => x"00", -- $0c22d
          49710 => x"00", -- $0c22e
          49711 => x"00", -- $0c22f
          49712 => x"00", -- $0c230
          49713 => x"00", -- $0c231
          49714 => x"00", -- $0c232
          49715 => x"00", -- $0c233
          49716 => x"00", -- $0c234
          49717 => x"00", -- $0c235
          49718 => x"00", -- $0c236
          49719 => x"00", -- $0c237
          49720 => x"00", -- $0c238
          49721 => x"00", -- $0c239
          49722 => x"00", -- $0c23a
          49723 => x"00", -- $0c23b
          49724 => x"00", -- $0c23c
          49725 => x"00", -- $0c23d
          49726 => x"00", -- $0c23e
          49727 => x"00", -- $0c23f
          49728 => x"00", -- $0c240
          49729 => x"00", -- $0c241
          49730 => x"00", -- $0c242
          49731 => x"00", -- $0c243
          49732 => x"00", -- $0c244
          49733 => x"00", -- $0c245
          49734 => x"00", -- $0c246
          49735 => x"00", -- $0c247
          49736 => x"00", -- $0c248
          49737 => x"00", -- $0c249
          49738 => x"00", -- $0c24a
          49739 => x"00", -- $0c24b
          49740 => x"00", -- $0c24c
          49741 => x"00", -- $0c24d
          49742 => x"00", -- $0c24e
          49743 => x"00", -- $0c24f
          49744 => x"00", -- $0c250
          49745 => x"00", -- $0c251
          49746 => x"00", -- $0c252
          49747 => x"00", -- $0c253
          49748 => x"00", -- $0c254
          49749 => x"00", -- $0c255
          49750 => x"00", -- $0c256
          49751 => x"00", -- $0c257
          49752 => x"00", -- $0c258
          49753 => x"00", -- $0c259
          49754 => x"00", -- $0c25a
          49755 => x"00", -- $0c25b
          49756 => x"00", -- $0c25c
          49757 => x"00", -- $0c25d
          49758 => x"00", -- $0c25e
          49759 => x"00", -- $0c25f
          49760 => x"00", -- $0c260
          49761 => x"00", -- $0c261
          49762 => x"00", -- $0c262
          49763 => x"00", -- $0c263
          49764 => x"00", -- $0c264
          49765 => x"00", -- $0c265
          49766 => x"00", -- $0c266
          49767 => x"00", -- $0c267
          49768 => x"00", -- $0c268
          49769 => x"00", -- $0c269
          49770 => x"00", -- $0c26a
          49771 => x"00", -- $0c26b
          49772 => x"00", -- $0c26c
          49773 => x"00", -- $0c26d
          49774 => x"00", -- $0c26e
          49775 => x"00", -- $0c26f
          49776 => x"00", -- $0c270
          49777 => x"00", -- $0c271
          49778 => x"00", -- $0c272
          49779 => x"00", -- $0c273
          49780 => x"00", -- $0c274
          49781 => x"00", -- $0c275
          49782 => x"00", -- $0c276
          49783 => x"00", -- $0c277
          49784 => x"00", -- $0c278
          49785 => x"00", -- $0c279
          49786 => x"00", -- $0c27a
          49787 => x"00", -- $0c27b
          49788 => x"00", -- $0c27c
          49789 => x"00", -- $0c27d
          49790 => x"00", -- $0c27e
          49791 => x"00", -- $0c27f
          49792 => x"00", -- $0c280
          49793 => x"00", -- $0c281
          49794 => x"00", -- $0c282
          49795 => x"00", -- $0c283
          49796 => x"00", -- $0c284
          49797 => x"00", -- $0c285
          49798 => x"00", -- $0c286
          49799 => x"00", -- $0c287
          49800 => x"00", -- $0c288
          49801 => x"00", -- $0c289
          49802 => x"00", -- $0c28a
          49803 => x"00", -- $0c28b
          49804 => x"00", -- $0c28c
          49805 => x"00", -- $0c28d
          49806 => x"00", -- $0c28e
          49807 => x"00", -- $0c28f
          49808 => x"00", -- $0c290
          49809 => x"00", -- $0c291
          49810 => x"00", -- $0c292
          49811 => x"00", -- $0c293
          49812 => x"00", -- $0c294
          49813 => x"00", -- $0c295
          49814 => x"00", -- $0c296
          49815 => x"00", -- $0c297
          49816 => x"00", -- $0c298
          49817 => x"00", -- $0c299
          49818 => x"00", -- $0c29a
          49819 => x"00", -- $0c29b
          49820 => x"00", -- $0c29c
          49821 => x"00", -- $0c29d
          49822 => x"00", -- $0c29e
          49823 => x"00", -- $0c29f
          49824 => x"00", -- $0c2a0
          49825 => x"00", -- $0c2a1
          49826 => x"00", -- $0c2a2
          49827 => x"00", -- $0c2a3
          49828 => x"00", -- $0c2a4
          49829 => x"00", -- $0c2a5
          49830 => x"00", -- $0c2a6
          49831 => x"00", -- $0c2a7
          49832 => x"00", -- $0c2a8
          49833 => x"00", -- $0c2a9
          49834 => x"00", -- $0c2aa
          49835 => x"00", -- $0c2ab
          49836 => x"00", -- $0c2ac
          49837 => x"00", -- $0c2ad
          49838 => x"00", -- $0c2ae
          49839 => x"00", -- $0c2af
          49840 => x"00", -- $0c2b0
          49841 => x"00", -- $0c2b1
          49842 => x"00", -- $0c2b2
          49843 => x"00", -- $0c2b3
          49844 => x"00", -- $0c2b4
          49845 => x"00", -- $0c2b5
          49846 => x"00", -- $0c2b6
          49847 => x"00", -- $0c2b7
          49848 => x"00", -- $0c2b8
          49849 => x"00", -- $0c2b9
          49850 => x"00", -- $0c2ba
          49851 => x"00", -- $0c2bb
          49852 => x"00", -- $0c2bc
          49853 => x"00", -- $0c2bd
          49854 => x"00", -- $0c2be
          49855 => x"00", -- $0c2bf
          49856 => x"00", -- $0c2c0
          49857 => x"00", -- $0c2c1
          49858 => x"00", -- $0c2c2
          49859 => x"00", -- $0c2c3
          49860 => x"00", -- $0c2c4
          49861 => x"00", -- $0c2c5
          49862 => x"00", -- $0c2c6
          49863 => x"00", -- $0c2c7
          49864 => x"00", -- $0c2c8
          49865 => x"00", -- $0c2c9
          49866 => x"00", -- $0c2ca
          49867 => x"00", -- $0c2cb
          49868 => x"00", -- $0c2cc
          49869 => x"00", -- $0c2cd
          49870 => x"00", -- $0c2ce
          49871 => x"00", -- $0c2cf
          49872 => x"00", -- $0c2d0
          49873 => x"00", -- $0c2d1
          49874 => x"00", -- $0c2d2
          49875 => x"00", -- $0c2d3
          49876 => x"00", -- $0c2d4
          49877 => x"00", -- $0c2d5
          49878 => x"00", -- $0c2d6
          49879 => x"00", -- $0c2d7
          49880 => x"00", -- $0c2d8
          49881 => x"00", -- $0c2d9
          49882 => x"00", -- $0c2da
          49883 => x"00", -- $0c2db
          49884 => x"00", -- $0c2dc
          49885 => x"00", -- $0c2dd
          49886 => x"00", -- $0c2de
          49887 => x"00", -- $0c2df
          49888 => x"00", -- $0c2e0
          49889 => x"00", -- $0c2e1
          49890 => x"00", -- $0c2e2
          49891 => x"00", -- $0c2e3
          49892 => x"00", -- $0c2e4
          49893 => x"00", -- $0c2e5
          49894 => x"00", -- $0c2e6
          49895 => x"00", -- $0c2e7
          49896 => x"00", -- $0c2e8
          49897 => x"00", -- $0c2e9
          49898 => x"00", -- $0c2ea
          49899 => x"00", -- $0c2eb
          49900 => x"00", -- $0c2ec
          49901 => x"00", -- $0c2ed
          49902 => x"00", -- $0c2ee
          49903 => x"00", -- $0c2ef
          49904 => x"00", -- $0c2f0
          49905 => x"00", -- $0c2f1
          49906 => x"00", -- $0c2f2
          49907 => x"00", -- $0c2f3
          49908 => x"00", -- $0c2f4
          49909 => x"00", -- $0c2f5
          49910 => x"00", -- $0c2f6
          49911 => x"00", -- $0c2f7
          49912 => x"00", -- $0c2f8
          49913 => x"00", -- $0c2f9
          49914 => x"00", -- $0c2fa
          49915 => x"00", -- $0c2fb
          49916 => x"00", -- $0c2fc
          49917 => x"00", -- $0c2fd
          49918 => x"00", -- $0c2fe
          49919 => x"00", -- $0c2ff
          49920 => x"00", -- $0c300
          49921 => x"00", -- $0c301
          49922 => x"00", -- $0c302
          49923 => x"00", -- $0c303
          49924 => x"00", -- $0c304
          49925 => x"00", -- $0c305
          49926 => x"00", -- $0c306
          49927 => x"00", -- $0c307
          49928 => x"00", -- $0c308
          49929 => x"00", -- $0c309
          49930 => x"00", -- $0c30a
          49931 => x"00", -- $0c30b
          49932 => x"00", -- $0c30c
          49933 => x"00", -- $0c30d
          49934 => x"00", -- $0c30e
          49935 => x"00", -- $0c30f
          49936 => x"00", -- $0c310
          49937 => x"00", -- $0c311
          49938 => x"00", -- $0c312
          49939 => x"00", -- $0c313
          49940 => x"00", -- $0c314
          49941 => x"00", -- $0c315
          49942 => x"00", -- $0c316
          49943 => x"00", -- $0c317
          49944 => x"00", -- $0c318
          49945 => x"00", -- $0c319
          49946 => x"00", -- $0c31a
          49947 => x"00", -- $0c31b
          49948 => x"00", -- $0c31c
          49949 => x"00", -- $0c31d
          49950 => x"00", -- $0c31e
          49951 => x"00", -- $0c31f
          49952 => x"00", -- $0c320
          49953 => x"00", -- $0c321
          49954 => x"00", -- $0c322
          49955 => x"00", -- $0c323
          49956 => x"00", -- $0c324
          49957 => x"00", -- $0c325
          49958 => x"00", -- $0c326
          49959 => x"00", -- $0c327
          49960 => x"00", -- $0c328
          49961 => x"00", -- $0c329
          49962 => x"00", -- $0c32a
          49963 => x"00", -- $0c32b
          49964 => x"00", -- $0c32c
          49965 => x"00", -- $0c32d
          49966 => x"00", -- $0c32e
          49967 => x"00", -- $0c32f
          49968 => x"00", -- $0c330
          49969 => x"00", -- $0c331
          49970 => x"00", -- $0c332
          49971 => x"00", -- $0c333
          49972 => x"00", -- $0c334
          49973 => x"00", -- $0c335
          49974 => x"00", -- $0c336
          49975 => x"00", -- $0c337
          49976 => x"00", -- $0c338
          49977 => x"00", -- $0c339
          49978 => x"00", -- $0c33a
          49979 => x"00", -- $0c33b
          49980 => x"00", -- $0c33c
          49981 => x"00", -- $0c33d
          49982 => x"00", -- $0c33e
          49983 => x"00", -- $0c33f
          49984 => x"00", -- $0c340
          49985 => x"00", -- $0c341
          49986 => x"00", -- $0c342
          49987 => x"00", -- $0c343
          49988 => x"00", -- $0c344
          49989 => x"00", -- $0c345
          49990 => x"00", -- $0c346
          49991 => x"00", -- $0c347
          49992 => x"00", -- $0c348
          49993 => x"00", -- $0c349
          49994 => x"00", -- $0c34a
          49995 => x"00", -- $0c34b
          49996 => x"00", -- $0c34c
          49997 => x"00", -- $0c34d
          49998 => x"00", -- $0c34e
          49999 => x"00", -- $0c34f
          50000 => x"00", -- $0c350
          50001 => x"00", -- $0c351
          50002 => x"00", -- $0c352
          50003 => x"00", -- $0c353
          50004 => x"00", -- $0c354
          50005 => x"00", -- $0c355
          50006 => x"00", -- $0c356
          50007 => x"00", -- $0c357
          50008 => x"00", -- $0c358
          50009 => x"00", -- $0c359
          50010 => x"00", -- $0c35a
          50011 => x"00", -- $0c35b
          50012 => x"00", -- $0c35c
          50013 => x"00", -- $0c35d
          50014 => x"00", -- $0c35e
          50015 => x"00", -- $0c35f
          50016 => x"00", -- $0c360
          50017 => x"00", -- $0c361
          50018 => x"00", -- $0c362
          50019 => x"00", -- $0c363
          50020 => x"00", -- $0c364
          50021 => x"00", -- $0c365
          50022 => x"00", -- $0c366
          50023 => x"00", -- $0c367
          50024 => x"00", -- $0c368
          50025 => x"00", -- $0c369
          50026 => x"00", -- $0c36a
          50027 => x"00", -- $0c36b
          50028 => x"00", -- $0c36c
          50029 => x"00", -- $0c36d
          50030 => x"00", -- $0c36e
          50031 => x"00", -- $0c36f
          50032 => x"00", -- $0c370
          50033 => x"00", -- $0c371
          50034 => x"00", -- $0c372
          50035 => x"00", -- $0c373
          50036 => x"00", -- $0c374
          50037 => x"00", -- $0c375
          50038 => x"00", -- $0c376
          50039 => x"00", -- $0c377
          50040 => x"00", -- $0c378
          50041 => x"00", -- $0c379
          50042 => x"00", -- $0c37a
          50043 => x"00", -- $0c37b
          50044 => x"00", -- $0c37c
          50045 => x"00", -- $0c37d
          50046 => x"00", -- $0c37e
          50047 => x"00", -- $0c37f
          50048 => x"00", -- $0c380
          50049 => x"00", -- $0c381
          50050 => x"00", -- $0c382
          50051 => x"00", -- $0c383
          50052 => x"00", -- $0c384
          50053 => x"00", -- $0c385
          50054 => x"00", -- $0c386
          50055 => x"00", -- $0c387
          50056 => x"00", -- $0c388
          50057 => x"00", -- $0c389
          50058 => x"00", -- $0c38a
          50059 => x"00", -- $0c38b
          50060 => x"00", -- $0c38c
          50061 => x"00", -- $0c38d
          50062 => x"00", -- $0c38e
          50063 => x"00", -- $0c38f
          50064 => x"00", -- $0c390
          50065 => x"00", -- $0c391
          50066 => x"00", -- $0c392
          50067 => x"00", -- $0c393
          50068 => x"00", -- $0c394
          50069 => x"00", -- $0c395
          50070 => x"00", -- $0c396
          50071 => x"00", -- $0c397
          50072 => x"00", -- $0c398
          50073 => x"00", -- $0c399
          50074 => x"00", -- $0c39a
          50075 => x"00", -- $0c39b
          50076 => x"00", -- $0c39c
          50077 => x"00", -- $0c39d
          50078 => x"00", -- $0c39e
          50079 => x"00", -- $0c39f
          50080 => x"00", -- $0c3a0
          50081 => x"00", -- $0c3a1
          50082 => x"00", -- $0c3a2
          50083 => x"00", -- $0c3a3
          50084 => x"00", -- $0c3a4
          50085 => x"00", -- $0c3a5
          50086 => x"00", -- $0c3a6
          50087 => x"00", -- $0c3a7
          50088 => x"00", -- $0c3a8
          50089 => x"00", -- $0c3a9
          50090 => x"00", -- $0c3aa
          50091 => x"00", -- $0c3ab
          50092 => x"00", -- $0c3ac
          50093 => x"00", -- $0c3ad
          50094 => x"00", -- $0c3ae
          50095 => x"00", -- $0c3af
          50096 => x"00", -- $0c3b0
          50097 => x"00", -- $0c3b1
          50098 => x"00", -- $0c3b2
          50099 => x"00", -- $0c3b3
          50100 => x"00", -- $0c3b4
          50101 => x"00", -- $0c3b5
          50102 => x"00", -- $0c3b6
          50103 => x"00", -- $0c3b7
          50104 => x"00", -- $0c3b8
          50105 => x"00", -- $0c3b9
          50106 => x"00", -- $0c3ba
          50107 => x"00", -- $0c3bb
          50108 => x"00", -- $0c3bc
          50109 => x"00", -- $0c3bd
          50110 => x"00", -- $0c3be
          50111 => x"00", -- $0c3bf
          50112 => x"00", -- $0c3c0
          50113 => x"00", -- $0c3c1
          50114 => x"00", -- $0c3c2
          50115 => x"00", -- $0c3c3
          50116 => x"00", -- $0c3c4
          50117 => x"00", -- $0c3c5
          50118 => x"00", -- $0c3c6
          50119 => x"00", -- $0c3c7
          50120 => x"00", -- $0c3c8
          50121 => x"00", -- $0c3c9
          50122 => x"00", -- $0c3ca
          50123 => x"00", -- $0c3cb
          50124 => x"00", -- $0c3cc
          50125 => x"00", -- $0c3cd
          50126 => x"00", -- $0c3ce
          50127 => x"00", -- $0c3cf
          50128 => x"00", -- $0c3d0
          50129 => x"00", -- $0c3d1
          50130 => x"00", -- $0c3d2
          50131 => x"00", -- $0c3d3
          50132 => x"00", -- $0c3d4
          50133 => x"00", -- $0c3d5
          50134 => x"00", -- $0c3d6
          50135 => x"00", -- $0c3d7
          50136 => x"00", -- $0c3d8
          50137 => x"00", -- $0c3d9
          50138 => x"00", -- $0c3da
          50139 => x"00", -- $0c3db
          50140 => x"00", -- $0c3dc
          50141 => x"00", -- $0c3dd
          50142 => x"00", -- $0c3de
          50143 => x"00", -- $0c3df
          50144 => x"00", -- $0c3e0
          50145 => x"00", -- $0c3e1
          50146 => x"00", -- $0c3e2
          50147 => x"00", -- $0c3e3
          50148 => x"00", -- $0c3e4
          50149 => x"00", -- $0c3e5
          50150 => x"00", -- $0c3e6
          50151 => x"00", -- $0c3e7
          50152 => x"00", -- $0c3e8
          50153 => x"00", -- $0c3e9
          50154 => x"00", -- $0c3ea
          50155 => x"00", -- $0c3eb
          50156 => x"00", -- $0c3ec
          50157 => x"00", -- $0c3ed
          50158 => x"00", -- $0c3ee
          50159 => x"00", -- $0c3ef
          50160 => x"00", -- $0c3f0
          50161 => x"00", -- $0c3f1
          50162 => x"00", -- $0c3f2
          50163 => x"00", -- $0c3f3
          50164 => x"00", -- $0c3f4
          50165 => x"00", -- $0c3f5
          50166 => x"00", -- $0c3f6
          50167 => x"00", -- $0c3f7
          50168 => x"00", -- $0c3f8
          50169 => x"00", -- $0c3f9
          50170 => x"00", -- $0c3fa
          50171 => x"00", -- $0c3fb
          50172 => x"00", -- $0c3fc
          50173 => x"00", -- $0c3fd
          50174 => x"00", -- $0c3fe
          50175 => x"00", -- $0c3ff
          50176 => x"00", -- $0c400
          50177 => x"00", -- $0c401
          50178 => x"00", -- $0c402
          50179 => x"00", -- $0c403
          50180 => x"00", -- $0c404
          50181 => x"00", -- $0c405
          50182 => x"00", -- $0c406
          50183 => x"00", -- $0c407
          50184 => x"00", -- $0c408
          50185 => x"00", -- $0c409
          50186 => x"00", -- $0c40a
          50187 => x"00", -- $0c40b
          50188 => x"00", -- $0c40c
          50189 => x"00", -- $0c40d
          50190 => x"00", -- $0c40e
          50191 => x"00", -- $0c40f
          50192 => x"00", -- $0c410
          50193 => x"00", -- $0c411
          50194 => x"00", -- $0c412
          50195 => x"00", -- $0c413
          50196 => x"00", -- $0c414
          50197 => x"00", -- $0c415
          50198 => x"00", -- $0c416
          50199 => x"00", -- $0c417
          50200 => x"00", -- $0c418
          50201 => x"00", -- $0c419
          50202 => x"00", -- $0c41a
          50203 => x"00", -- $0c41b
          50204 => x"00", -- $0c41c
          50205 => x"00", -- $0c41d
          50206 => x"00", -- $0c41e
          50207 => x"00", -- $0c41f
          50208 => x"00", -- $0c420
          50209 => x"00", -- $0c421
          50210 => x"00", -- $0c422
          50211 => x"00", -- $0c423
          50212 => x"00", -- $0c424
          50213 => x"00", -- $0c425
          50214 => x"00", -- $0c426
          50215 => x"00", -- $0c427
          50216 => x"00", -- $0c428
          50217 => x"00", -- $0c429
          50218 => x"00", -- $0c42a
          50219 => x"00", -- $0c42b
          50220 => x"00", -- $0c42c
          50221 => x"00", -- $0c42d
          50222 => x"00", -- $0c42e
          50223 => x"00", -- $0c42f
          50224 => x"00", -- $0c430
          50225 => x"00", -- $0c431
          50226 => x"00", -- $0c432
          50227 => x"00", -- $0c433
          50228 => x"00", -- $0c434
          50229 => x"00", -- $0c435
          50230 => x"00", -- $0c436
          50231 => x"00", -- $0c437
          50232 => x"00", -- $0c438
          50233 => x"00", -- $0c439
          50234 => x"00", -- $0c43a
          50235 => x"00", -- $0c43b
          50236 => x"00", -- $0c43c
          50237 => x"00", -- $0c43d
          50238 => x"00", -- $0c43e
          50239 => x"00", -- $0c43f
          50240 => x"00", -- $0c440
          50241 => x"00", -- $0c441
          50242 => x"00", -- $0c442
          50243 => x"00", -- $0c443
          50244 => x"00", -- $0c444
          50245 => x"00", -- $0c445
          50246 => x"00", -- $0c446
          50247 => x"00", -- $0c447
          50248 => x"00", -- $0c448
          50249 => x"00", -- $0c449
          50250 => x"00", -- $0c44a
          50251 => x"00", -- $0c44b
          50252 => x"00", -- $0c44c
          50253 => x"00", -- $0c44d
          50254 => x"00", -- $0c44e
          50255 => x"00", -- $0c44f
          50256 => x"00", -- $0c450
          50257 => x"00", -- $0c451
          50258 => x"00", -- $0c452
          50259 => x"00", -- $0c453
          50260 => x"00", -- $0c454
          50261 => x"00", -- $0c455
          50262 => x"00", -- $0c456
          50263 => x"00", -- $0c457
          50264 => x"00", -- $0c458
          50265 => x"00", -- $0c459
          50266 => x"00", -- $0c45a
          50267 => x"00", -- $0c45b
          50268 => x"00", -- $0c45c
          50269 => x"00", -- $0c45d
          50270 => x"00", -- $0c45e
          50271 => x"00", -- $0c45f
          50272 => x"00", -- $0c460
          50273 => x"00", -- $0c461
          50274 => x"00", -- $0c462
          50275 => x"00", -- $0c463
          50276 => x"00", -- $0c464
          50277 => x"00", -- $0c465
          50278 => x"00", -- $0c466
          50279 => x"00", -- $0c467
          50280 => x"00", -- $0c468
          50281 => x"00", -- $0c469
          50282 => x"00", -- $0c46a
          50283 => x"00", -- $0c46b
          50284 => x"00", -- $0c46c
          50285 => x"00", -- $0c46d
          50286 => x"00", -- $0c46e
          50287 => x"00", -- $0c46f
          50288 => x"00", -- $0c470
          50289 => x"00", -- $0c471
          50290 => x"00", -- $0c472
          50291 => x"00", -- $0c473
          50292 => x"00", -- $0c474
          50293 => x"00", -- $0c475
          50294 => x"00", -- $0c476
          50295 => x"00", -- $0c477
          50296 => x"00", -- $0c478
          50297 => x"00", -- $0c479
          50298 => x"00", -- $0c47a
          50299 => x"00", -- $0c47b
          50300 => x"00", -- $0c47c
          50301 => x"00", -- $0c47d
          50302 => x"00", -- $0c47e
          50303 => x"00", -- $0c47f
          50304 => x"00", -- $0c480
          50305 => x"00", -- $0c481
          50306 => x"00", -- $0c482
          50307 => x"00", -- $0c483
          50308 => x"00", -- $0c484
          50309 => x"00", -- $0c485
          50310 => x"00", -- $0c486
          50311 => x"00", -- $0c487
          50312 => x"00", -- $0c488
          50313 => x"00", -- $0c489
          50314 => x"00", -- $0c48a
          50315 => x"00", -- $0c48b
          50316 => x"00", -- $0c48c
          50317 => x"00", -- $0c48d
          50318 => x"00", -- $0c48e
          50319 => x"00", -- $0c48f
          50320 => x"00", -- $0c490
          50321 => x"00", -- $0c491
          50322 => x"00", -- $0c492
          50323 => x"00", -- $0c493
          50324 => x"00", -- $0c494
          50325 => x"00", -- $0c495
          50326 => x"00", -- $0c496
          50327 => x"00", -- $0c497
          50328 => x"00", -- $0c498
          50329 => x"00", -- $0c499
          50330 => x"00", -- $0c49a
          50331 => x"00", -- $0c49b
          50332 => x"00", -- $0c49c
          50333 => x"00", -- $0c49d
          50334 => x"00", -- $0c49e
          50335 => x"00", -- $0c49f
          50336 => x"00", -- $0c4a0
          50337 => x"00", -- $0c4a1
          50338 => x"00", -- $0c4a2
          50339 => x"00", -- $0c4a3
          50340 => x"00", -- $0c4a4
          50341 => x"00", -- $0c4a5
          50342 => x"00", -- $0c4a6
          50343 => x"00", -- $0c4a7
          50344 => x"00", -- $0c4a8
          50345 => x"00", -- $0c4a9
          50346 => x"00", -- $0c4aa
          50347 => x"00", -- $0c4ab
          50348 => x"00", -- $0c4ac
          50349 => x"00", -- $0c4ad
          50350 => x"00", -- $0c4ae
          50351 => x"00", -- $0c4af
          50352 => x"00", -- $0c4b0
          50353 => x"00", -- $0c4b1
          50354 => x"00", -- $0c4b2
          50355 => x"00", -- $0c4b3
          50356 => x"00", -- $0c4b4
          50357 => x"00", -- $0c4b5
          50358 => x"00", -- $0c4b6
          50359 => x"00", -- $0c4b7
          50360 => x"00", -- $0c4b8
          50361 => x"00", -- $0c4b9
          50362 => x"00", -- $0c4ba
          50363 => x"00", -- $0c4bb
          50364 => x"00", -- $0c4bc
          50365 => x"00", -- $0c4bd
          50366 => x"00", -- $0c4be
          50367 => x"00", -- $0c4bf
          50368 => x"00", -- $0c4c0
          50369 => x"00", -- $0c4c1
          50370 => x"00", -- $0c4c2
          50371 => x"00", -- $0c4c3
          50372 => x"00", -- $0c4c4
          50373 => x"00", -- $0c4c5
          50374 => x"00", -- $0c4c6
          50375 => x"00", -- $0c4c7
          50376 => x"00", -- $0c4c8
          50377 => x"00", -- $0c4c9
          50378 => x"00", -- $0c4ca
          50379 => x"00", -- $0c4cb
          50380 => x"00", -- $0c4cc
          50381 => x"00", -- $0c4cd
          50382 => x"00", -- $0c4ce
          50383 => x"00", -- $0c4cf
          50384 => x"00", -- $0c4d0
          50385 => x"00", -- $0c4d1
          50386 => x"00", -- $0c4d2
          50387 => x"00", -- $0c4d3
          50388 => x"00", -- $0c4d4
          50389 => x"00", -- $0c4d5
          50390 => x"00", -- $0c4d6
          50391 => x"00", -- $0c4d7
          50392 => x"00", -- $0c4d8
          50393 => x"00", -- $0c4d9
          50394 => x"00", -- $0c4da
          50395 => x"00", -- $0c4db
          50396 => x"00", -- $0c4dc
          50397 => x"00", -- $0c4dd
          50398 => x"00", -- $0c4de
          50399 => x"00", -- $0c4df
          50400 => x"00", -- $0c4e0
          50401 => x"00", -- $0c4e1
          50402 => x"00", -- $0c4e2
          50403 => x"00", -- $0c4e3
          50404 => x"00", -- $0c4e4
          50405 => x"00", -- $0c4e5
          50406 => x"00", -- $0c4e6
          50407 => x"00", -- $0c4e7
          50408 => x"00", -- $0c4e8
          50409 => x"00", -- $0c4e9
          50410 => x"00", -- $0c4ea
          50411 => x"00", -- $0c4eb
          50412 => x"00", -- $0c4ec
          50413 => x"00", -- $0c4ed
          50414 => x"00", -- $0c4ee
          50415 => x"00", -- $0c4ef
          50416 => x"00", -- $0c4f0
          50417 => x"00", -- $0c4f1
          50418 => x"00", -- $0c4f2
          50419 => x"00", -- $0c4f3
          50420 => x"00", -- $0c4f4
          50421 => x"00", -- $0c4f5
          50422 => x"00", -- $0c4f6
          50423 => x"00", -- $0c4f7
          50424 => x"00", -- $0c4f8
          50425 => x"00", -- $0c4f9
          50426 => x"00", -- $0c4fa
          50427 => x"00", -- $0c4fb
          50428 => x"00", -- $0c4fc
          50429 => x"00", -- $0c4fd
          50430 => x"00", -- $0c4fe
          50431 => x"00", -- $0c4ff
          50432 => x"00", -- $0c500
          50433 => x"00", -- $0c501
          50434 => x"00", -- $0c502
          50435 => x"00", -- $0c503
          50436 => x"00", -- $0c504
          50437 => x"00", -- $0c505
          50438 => x"00", -- $0c506
          50439 => x"00", -- $0c507
          50440 => x"00", -- $0c508
          50441 => x"00", -- $0c509
          50442 => x"00", -- $0c50a
          50443 => x"00", -- $0c50b
          50444 => x"00", -- $0c50c
          50445 => x"00", -- $0c50d
          50446 => x"00", -- $0c50e
          50447 => x"00", -- $0c50f
          50448 => x"00", -- $0c510
          50449 => x"00", -- $0c511
          50450 => x"00", -- $0c512
          50451 => x"00", -- $0c513
          50452 => x"00", -- $0c514
          50453 => x"00", -- $0c515
          50454 => x"00", -- $0c516
          50455 => x"00", -- $0c517
          50456 => x"00", -- $0c518
          50457 => x"00", -- $0c519
          50458 => x"00", -- $0c51a
          50459 => x"00", -- $0c51b
          50460 => x"00", -- $0c51c
          50461 => x"00", -- $0c51d
          50462 => x"00", -- $0c51e
          50463 => x"00", -- $0c51f
          50464 => x"00", -- $0c520
          50465 => x"00", -- $0c521
          50466 => x"00", -- $0c522
          50467 => x"00", -- $0c523
          50468 => x"00", -- $0c524
          50469 => x"00", -- $0c525
          50470 => x"00", -- $0c526
          50471 => x"00", -- $0c527
          50472 => x"00", -- $0c528
          50473 => x"00", -- $0c529
          50474 => x"00", -- $0c52a
          50475 => x"00", -- $0c52b
          50476 => x"00", -- $0c52c
          50477 => x"00", -- $0c52d
          50478 => x"00", -- $0c52e
          50479 => x"00", -- $0c52f
          50480 => x"00", -- $0c530
          50481 => x"00", -- $0c531
          50482 => x"00", -- $0c532
          50483 => x"00", -- $0c533
          50484 => x"00", -- $0c534
          50485 => x"00", -- $0c535
          50486 => x"00", -- $0c536
          50487 => x"00", -- $0c537
          50488 => x"00", -- $0c538
          50489 => x"00", -- $0c539
          50490 => x"00", -- $0c53a
          50491 => x"00", -- $0c53b
          50492 => x"00", -- $0c53c
          50493 => x"00", -- $0c53d
          50494 => x"00", -- $0c53e
          50495 => x"00", -- $0c53f
          50496 => x"00", -- $0c540
          50497 => x"00", -- $0c541
          50498 => x"00", -- $0c542
          50499 => x"00", -- $0c543
          50500 => x"00", -- $0c544
          50501 => x"00", -- $0c545
          50502 => x"00", -- $0c546
          50503 => x"00", -- $0c547
          50504 => x"00", -- $0c548
          50505 => x"00", -- $0c549
          50506 => x"00", -- $0c54a
          50507 => x"00", -- $0c54b
          50508 => x"00", -- $0c54c
          50509 => x"00", -- $0c54d
          50510 => x"00", -- $0c54e
          50511 => x"00", -- $0c54f
          50512 => x"00", -- $0c550
          50513 => x"00", -- $0c551
          50514 => x"00", -- $0c552
          50515 => x"00", -- $0c553
          50516 => x"00", -- $0c554
          50517 => x"00", -- $0c555
          50518 => x"00", -- $0c556
          50519 => x"00", -- $0c557
          50520 => x"00", -- $0c558
          50521 => x"00", -- $0c559
          50522 => x"00", -- $0c55a
          50523 => x"00", -- $0c55b
          50524 => x"00", -- $0c55c
          50525 => x"00", -- $0c55d
          50526 => x"00", -- $0c55e
          50527 => x"00", -- $0c55f
          50528 => x"00", -- $0c560
          50529 => x"00", -- $0c561
          50530 => x"00", -- $0c562
          50531 => x"00", -- $0c563
          50532 => x"00", -- $0c564
          50533 => x"00", -- $0c565
          50534 => x"00", -- $0c566
          50535 => x"00", -- $0c567
          50536 => x"00", -- $0c568
          50537 => x"00", -- $0c569
          50538 => x"00", -- $0c56a
          50539 => x"00", -- $0c56b
          50540 => x"00", -- $0c56c
          50541 => x"00", -- $0c56d
          50542 => x"00", -- $0c56e
          50543 => x"00", -- $0c56f
          50544 => x"00", -- $0c570
          50545 => x"00", -- $0c571
          50546 => x"00", -- $0c572
          50547 => x"00", -- $0c573
          50548 => x"00", -- $0c574
          50549 => x"00", -- $0c575
          50550 => x"00", -- $0c576
          50551 => x"00", -- $0c577
          50552 => x"00", -- $0c578
          50553 => x"00", -- $0c579
          50554 => x"00", -- $0c57a
          50555 => x"00", -- $0c57b
          50556 => x"00", -- $0c57c
          50557 => x"00", -- $0c57d
          50558 => x"00", -- $0c57e
          50559 => x"00", -- $0c57f
          50560 => x"00", -- $0c580
          50561 => x"00", -- $0c581
          50562 => x"00", -- $0c582
          50563 => x"00", -- $0c583
          50564 => x"00", -- $0c584
          50565 => x"00", -- $0c585
          50566 => x"00", -- $0c586
          50567 => x"00", -- $0c587
          50568 => x"00", -- $0c588
          50569 => x"00", -- $0c589
          50570 => x"00", -- $0c58a
          50571 => x"00", -- $0c58b
          50572 => x"00", -- $0c58c
          50573 => x"00", -- $0c58d
          50574 => x"00", -- $0c58e
          50575 => x"00", -- $0c58f
          50576 => x"00", -- $0c590
          50577 => x"00", -- $0c591
          50578 => x"00", -- $0c592
          50579 => x"00", -- $0c593
          50580 => x"00", -- $0c594
          50581 => x"00", -- $0c595
          50582 => x"00", -- $0c596
          50583 => x"00", -- $0c597
          50584 => x"00", -- $0c598
          50585 => x"00", -- $0c599
          50586 => x"00", -- $0c59a
          50587 => x"00", -- $0c59b
          50588 => x"00", -- $0c59c
          50589 => x"00", -- $0c59d
          50590 => x"00", -- $0c59e
          50591 => x"00", -- $0c59f
          50592 => x"00", -- $0c5a0
          50593 => x"00", -- $0c5a1
          50594 => x"00", -- $0c5a2
          50595 => x"00", -- $0c5a3
          50596 => x"00", -- $0c5a4
          50597 => x"00", -- $0c5a5
          50598 => x"00", -- $0c5a6
          50599 => x"00", -- $0c5a7
          50600 => x"00", -- $0c5a8
          50601 => x"00", -- $0c5a9
          50602 => x"00", -- $0c5aa
          50603 => x"00", -- $0c5ab
          50604 => x"00", -- $0c5ac
          50605 => x"00", -- $0c5ad
          50606 => x"00", -- $0c5ae
          50607 => x"00", -- $0c5af
          50608 => x"00", -- $0c5b0
          50609 => x"00", -- $0c5b1
          50610 => x"00", -- $0c5b2
          50611 => x"00", -- $0c5b3
          50612 => x"00", -- $0c5b4
          50613 => x"00", -- $0c5b5
          50614 => x"00", -- $0c5b6
          50615 => x"00", -- $0c5b7
          50616 => x"00", -- $0c5b8
          50617 => x"00", -- $0c5b9
          50618 => x"00", -- $0c5ba
          50619 => x"00", -- $0c5bb
          50620 => x"00", -- $0c5bc
          50621 => x"00", -- $0c5bd
          50622 => x"00", -- $0c5be
          50623 => x"00", -- $0c5bf
          50624 => x"00", -- $0c5c0
          50625 => x"00", -- $0c5c1
          50626 => x"00", -- $0c5c2
          50627 => x"00", -- $0c5c3
          50628 => x"00", -- $0c5c4
          50629 => x"00", -- $0c5c5
          50630 => x"00", -- $0c5c6
          50631 => x"00", -- $0c5c7
          50632 => x"00", -- $0c5c8
          50633 => x"00", -- $0c5c9
          50634 => x"00", -- $0c5ca
          50635 => x"00", -- $0c5cb
          50636 => x"00", -- $0c5cc
          50637 => x"00", -- $0c5cd
          50638 => x"00", -- $0c5ce
          50639 => x"00", -- $0c5cf
          50640 => x"00", -- $0c5d0
          50641 => x"00", -- $0c5d1
          50642 => x"00", -- $0c5d2
          50643 => x"00", -- $0c5d3
          50644 => x"00", -- $0c5d4
          50645 => x"00", -- $0c5d5
          50646 => x"00", -- $0c5d6
          50647 => x"00", -- $0c5d7
          50648 => x"00", -- $0c5d8
          50649 => x"00", -- $0c5d9
          50650 => x"00", -- $0c5da
          50651 => x"00", -- $0c5db
          50652 => x"00", -- $0c5dc
          50653 => x"00", -- $0c5dd
          50654 => x"00", -- $0c5de
          50655 => x"00", -- $0c5df
          50656 => x"00", -- $0c5e0
          50657 => x"00", -- $0c5e1
          50658 => x"00", -- $0c5e2
          50659 => x"00", -- $0c5e3
          50660 => x"00", -- $0c5e4
          50661 => x"00", -- $0c5e5
          50662 => x"00", -- $0c5e6
          50663 => x"00", -- $0c5e7
          50664 => x"00", -- $0c5e8
          50665 => x"00", -- $0c5e9
          50666 => x"00", -- $0c5ea
          50667 => x"00", -- $0c5eb
          50668 => x"00", -- $0c5ec
          50669 => x"00", -- $0c5ed
          50670 => x"00", -- $0c5ee
          50671 => x"00", -- $0c5ef
          50672 => x"00", -- $0c5f0
          50673 => x"00", -- $0c5f1
          50674 => x"00", -- $0c5f2
          50675 => x"00", -- $0c5f3
          50676 => x"00", -- $0c5f4
          50677 => x"00", -- $0c5f5
          50678 => x"00", -- $0c5f6
          50679 => x"00", -- $0c5f7
          50680 => x"00", -- $0c5f8
          50681 => x"00", -- $0c5f9
          50682 => x"00", -- $0c5fa
          50683 => x"00", -- $0c5fb
          50684 => x"00", -- $0c5fc
          50685 => x"00", -- $0c5fd
          50686 => x"00", -- $0c5fe
          50687 => x"00", -- $0c5ff
          50688 => x"00", -- $0c600
          50689 => x"00", -- $0c601
          50690 => x"00", -- $0c602
          50691 => x"00", -- $0c603
          50692 => x"00", -- $0c604
          50693 => x"00", -- $0c605
          50694 => x"00", -- $0c606
          50695 => x"00", -- $0c607
          50696 => x"00", -- $0c608
          50697 => x"00", -- $0c609
          50698 => x"00", -- $0c60a
          50699 => x"00", -- $0c60b
          50700 => x"00", -- $0c60c
          50701 => x"00", -- $0c60d
          50702 => x"00", -- $0c60e
          50703 => x"00", -- $0c60f
          50704 => x"00", -- $0c610
          50705 => x"00", -- $0c611
          50706 => x"00", -- $0c612
          50707 => x"00", -- $0c613
          50708 => x"00", -- $0c614
          50709 => x"00", -- $0c615
          50710 => x"00", -- $0c616
          50711 => x"00", -- $0c617
          50712 => x"00", -- $0c618
          50713 => x"00", -- $0c619
          50714 => x"00", -- $0c61a
          50715 => x"00", -- $0c61b
          50716 => x"00", -- $0c61c
          50717 => x"00", -- $0c61d
          50718 => x"00", -- $0c61e
          50719 => x"00", -- $0c61f
          50720 => x"00", -- $0c620
          50721 => x"00", -- $0c621
          50722 => x"00", -- $0c622
          50723 => x"00", -- $0c623
          50724 => x"00", -- $0c624
          50725 => x"00", -- $0c625
          50726 => x"00", -- $0c626
          50727 => x"00", -- $0c627
          50728 => x"00", -- $0c628
          50729 => x"00", -- $0c629
          50730 => x"00", -- $0c62a
          50731 => x"00", -- $0c62b
          50732 => x"00", -- $0c62c
          50733 => x"00", -- $0c62d
          50734 => x"00", -- $0c62e
          50735 => x"00", -- $0c62f
          50736 => x"00", -- $0c630
          50737 => x"00", -- $0c631
          50738 => x"00", -- $0c632
          50739 => x"00", -- $0c633
          50740 => x"00", -- $0c634
          50741 => x"00", -- $0c635
          50742 => x"00", -- $0c636
          50743 => x"00", -- $0c637
          50744 => x"00", -- $0c638
          50745 => x"00", -- $0c639
          50746 => x"00", -- $0c63a
          50747 => x"00", -- $0c63b
          50748 => x"00", -- $0c63c
          50749 => x"00", -- $0c63d
          50750 => x"00", -- $0c63e
          50751 => x"00", -- $0c63f
          50752 => x"00", -- $0c640
          50753 => x"00", -- $0c641
          50754 => x"00", -- $0c642
          50755 => x"00", -- $0c643
          50756 => x"00", -- $0c644
          50757 => x"00", -- $0c645
          50758 => x"00", -- $0c646
          50759 => x"00", -- $0c647
          50760 => x"00", -- $0c648
          50761 => x"00", -- $0c649
          50762 => x"00", -- $0c64a
          50763 => x"00", -- $0c64b
          50764 => x"00", -- $0c64c
          50765 => x"00", -- $0c64d
          50766 => x"00", -- $0c64e
          50767 => x"00", -- $0c64f
          50768 => x"00", -- $0c650
          50769 => x"00", -- $0c651
          50770 => x"00", -- $0c652
          50771 => x"00", -- $0c653
          50772 => x"00", -- $0c654
          50773 => x"00", -- $0c655
          50774 => x"00", -- $0c656
          50775 => x"00", -- $0c657
          50776 => x"00", -- $0c658
          50777 => x"00", -- $0c659
          50778 => x"00", -- $0c65a
          50779 => x"00", -- $0c65b
          50780 => x"00", -- $0c65c
          50781 => x"00", -- $0c65d
          50782 => x"00", -- $0c65e
          50783 => x"00", -- $0c65f
          50784 => x"00", -- $0c660
          50785 => x"00", -- $0c661
          50786 => x"00", -- $0c662
          50787 => x"00", -- $0c663
          50788 => x"00", -- $0c664
          50789 => x"00", -- $0c665
          50790 => x"00", -- $0c666
          50791 => x"00", -- $0c667
          50792 => x"00", -- $0c668
          50793 => x"00", -- $0c669
          50794 => x"00", -- $0c66a
          50795 => x"00", -- $0c66b
          50796 => x"00", -- $0c66c
          50797 => x"00", -- $0c66d
          50798 => x"00", -- $0c66e
          50799 => x"00", -- $0c66f
          50800 => x"00", -- $0c670
          50801 => x"00", -- $0c671
          50802 => x"00", -- $0c672
          50803 => x"00", -- $0c673
          50804 => x"00", -- $0c674
          50805 => x"00", -- $0c675
          50806 => x"00", -- $0c676
          50807 => x"00", -- $0c677
          50808 => x"00", -- $0c678
          50809 => x"00", -- $0c679
          50810 => x"00", -- $0c67a
          50811 => x"00", -- $0c67b
          50812 => x"00", -- $0c67c
          50813 => x"00", -- $0c67d
          50814 => x"00", -- $0c67e
          50815 => x"00", -- $0c67f
          50816 => x"00", -- $0c680
          50817 => x"00", -- $0c681
          50818 => x"00", -- $0c682
          50819 => x"00", -- $0c683
          50820 => x"00", -- $0c684
          50821 => x"00", -- $0c685
          50822 => x"00", -- $0c686
          50823 => x"00", -- $0c687
          50824 => x"00", -- $0c688
          50825 => x"00", -- $0c689
          50826 => x"00", -- $0c68a
          50827 => x"00", -- $0c68b
          50828 => x"00", -- $0c68c
          50829 => x"00", -- $0c68d
          50830 => x"00", -- $0c68e
          50831 => x"00", -- $0c68f
          50832 => x"00", -- $0c690
          50833 => x"00", -- $0c691
          50834 => x"00", -- $0c692
          50835 => x"00", -- $0c693
          50836 => x"00", -- $0c694
          50837 => x"00", -- $0c695
          50838 => x"00", -- $0c696
          50839 => x"00", -- $0c697
          50840 => x"00", -- $0c698
          50841 => x"00", -- $0c699
          50842 => x"00", -- $0c69a
          50843 => x"00", -- $0c69b
          50844 => x"00", -- $0c69c
          50845 => x"00", -- $0c69d
          50846 => x"00", -- $0c69e
          50847 => x"00", -- $0c69f
          50848 => x"00", -- $0c6a0
          50849 => x"00", -- $0c6a1
          50850 => x"00", -- $0c6a2
          50851 => x"00", -- $0c6a3
          50852 => x"00", -- $0c6a4
          50853 => x"00", -- $0c6a5
          50854 => x"00", -- $0c6a6
          50855 => x"00", -- $0c6a7
          50856 => x"00", -- $0c6a8
          50857 => x"00", -- $0c6a9
          50858 => x"00", -- $0c6aa
          50859 => x"00", -- $0c6ab
          50860 => x"00", -- $0c6ac
          50861 => x"00", -- $0c6ad
          50862 => x"00", -- $0c6ae
          50863 => x"00", -- $0c6af
          50864 => x"00", -- $0c6b0
          50865 => x"00", -- $0c6b1
          50866 => x"00", -- $0c6b2
          50867 => x"00", -- $0c6b3
          50868 => x"00", -- $0c6b4
          50869 => x"00", -- $0c6b5
          50870 => x"00", -- $0c6b6
          50871 => x"00", -- $0c6b7
          50872 => x"00", -- $0c6b8
          50873 => x"00", -- $0c6b9
          50874 => x"00", -- $0c6ba
          50875 => x"00", -- $0c6bb
          50876 => x"00", -- $0c6bc
          50877 => x"00", -- $0c6bd
          50878 => x"00", -- $0c6be
          50879 => x"00", -- $0c6bf
          50880 => x"00", -- $0c6c0
          50881 => x"00", -- $0c6c1
          50882 => x"00", -- $0c6c2
          50883 => x"00", -- $0c6c3
          50884 => x"00", -- $0c6c4
          50885 => x"00", -- $0c6c5
          50886 => x"00", -- $0c6c6
          50887 => x"00", -- $0c6c7
          50888 => x"00", -- $0c6c8
          50889 => x"00", -- $0c6c9
          50890 => x"00", -- $0c6ca
          50891 => x"00", -- $0c6cb
          50892 => x"00", -- $0c6cc
          50893 => x"00", -- $0c6cd
          50894 => x"00", -- $0c6ce
          50895 => x"00", -- $0c6cf
          50896 => x"00", -- $0c6d0
          50897 => x"00", -- $0c6d1
          50898 => x"00", -- $0c6d2
          50899 => x"00", -- $0c6d3
          50900 => x"00", -- $0c6d4
          50901 => x"00", -- $0c6d5
          50902 => x"00", -- $0c6d6
          50903 => x"00", -- $0c6d7
          50904 => x"00", -- $0c6d8
          50905 => x"00", -- $0c6d9
          50906 => x"00", -- $0c6da
          50907 => x"00", -- $0c6db
          50908 => x"00", -- $0c6dc
          50909 => x"00", -- $0c6dd
          50910 => x"00", -- $0c6de
          50911 => x"00", -- $0c6df
          50912 => x"00", -- $0c6e0
          50913 => x"00", -- $0c6e1
          50914 => x"00", -- $0c6e2
          50915 => x"00", -- $0c6e3
          50916 => x"00", -- $0c6e4
          50917 => x"00", -- $0c6e5
          50918 => x"00", -- $0c6e6
          50919 => x"00", -- $0c6e7
          50920 => x"00", -- $0c6e8
          50921 => x"00", -- $0c6e9
          50922 => x"00", -- $0c6ea
          50923 => x"00", -- $0c6eb
          50924 => x"00", -- $0c6ec
          50925 => x"00", -- $0c6ed
          50926 => x"00", -- $0c6ee
          50927 => x"00", -- $0c6ef
          50928 => x"00", -- $0c6f0
          50929 => x"00", -- $0c6f1
          50930 => x"00", -- $0c6f2
          50931 => x"00", -- $0c6f3
          50932 => x"00", -- $0c6f4
          50933 => x"00", -- $0c6f5
          50934 => x"00", -- $0c6f6
          50935 => x"00", -- $0c6f7
          50936 => x"00", -- $0c6f8
          50937 => x"00", -- $0c6f9
          50938 => x"00", -- $0c6fa
          50939 => x"00", -- $0c6fb
          50940 => x"00", -- $0c6fc
          50941 => x"00", -- $0c6fd
          50942 => x"00", -- $0c6fe
          50943 => x"00", -- $0c6ff
          50944 => x"00", -- $0c700
          50945 => x"00", -- $0c701
          50946 => x"00", -- $0c702
          50947 => x"00", -- $0c703
          50948 => x"00", -- $0c704
          50949 => x"00", -- $0c705
          50950 => x"00", -- $0c706
          50951 => x"00", -- $0c707
          50952 => x"00", -- $0c708
          50953 => x"00", -- $0c709
          50954 => x"00", -- $0c70a
          50955 => x"00", -- $0c70b
          50956 => x"00", -- $0c70c
          50957 => x"00", -- $0c70d
          50958 => x"00", -- $0c70e
          50959 => x"00", -- $0c70f
          50960 => x"00", -- $0c710
          50961 => x"00", -- $0c711
          50962 => x"00", -- $0c712
          50963 => x"00", -- $0c713
          50964 => x"00", -- $0c714
          50965 => x"00", -- $0c715
          50966 => x"00", -- $0c716
          50967 => x"00", -- $0c717
          50968 => x"00", -- $0c718
          50969 => x"00", -- $0c719
          50970 => x"00", -- $0c71a
          50971 => x"00", -- $0c71b
          50972 => x"00", -- $0c71c
          50973 => x"00", -- $0c71d
          50974 => x"00", -- $0c71e
          50975 => x"00", -- $0c71f
          50976 => x"00", -- $0c720
          50977 => x"00", -- $0c721
          50978 => x"00", -- $0c722
          50979 => x"00", -- $0c723
          50980 => x"00", -- $0c724
          50981 => x"00", -- $0c725
          50982 => x"00", -- $0c726
          50983 => x"00", -- $0c727
          50984 => x"00", -- $0c728
          50985 => x"00", -- $0c729
          50986 => x"00", -- $0c72a
          50987 => x"00", -- $0c72b
          50988 => x"00", -- $0c72c
          50989 => x"00", -- $0c72d
          50990 => x"00", -- $0c72e
          50991 => x"00", -- $0c72f
          50992 => x"00", -- $0c730
          50993 => x"00", -- $0c731
          50994 => x"00", -- $0c732
          50995 => x"00", -- $0c733
          50996 => x"00", -- $0c734
          50997 => x"00", -- $0c735
          50998 => x"00", -- $0c736
          50999 => x"00", -- $0c737
          51000 => x"00", -- $0c738
          51001 => x"00", -- $0c739
          51002 => x"00", -- $0c73a
          51003 => x"00", -- $0c73b
          51004 => x"00", -- $0c73c
          51005 => x"00", -- $0c73d
          51006 => x"00", -- $0c73e
          51007 => x"00", -- $0c73f
          51008 => x"00", -- $0c740
          51009 => x"00", -- $0c741
          51010 => x"00", -- $0c742
          51011 => x"00", -- $0c743
          51012 => x"00", -- $0c744
          51013 => x"00", -- $0c745
          51014 => x"00", -- $0c746
          51015 => x"00", -- $0c747
          51016 => x"00", -- $0c748
          51017 => x"00", -- $0c749
          51018 => x"00", -- $0c74a
          51019 => x"00", -- $0c74b
          51020 => x"00", -- $0c74c
          51021 => x"00", -- $0c74d
          51022 => x"00", -- $0c74e
          51023 => x"00", -- $0c74f
          51024 => x"00", -- $0c750
          51025 => x"00", -- $0c751
          51026 => x"00", -- $0c752
          51027 => x"00", -- $0c753
          51028 => x"00", -- $0c754
          51029 => x"00", -- $0c755
          51030 => x"00", -- $0c756
          51031 => x"00", -- $0c757
          51032 => x"00", -- $0c758
          51033 => x"00", -- $0c759
          51034 => x"00", -- $0c75a
          51035 => x"00", -- $0c75b
          51036 => x"00", -- $0c75c
          51037 => x"00", -- $0c75d
          51038 => x"00", -- $0c75e
          51039 => x"00", -- $0c75f
          51040 => x"00", -- $0c760
          51041 => x"00", -- $0c761
          51042 => x"00", -- $0c762
          51043 => x"00", -- $0c763
          51044 => x"00", -- $0c764
          51045 => x"00", -- $0c765
          51046 => x"00", -- $0c766
          51047 => x"00", -- $0c767
          51048 => x"00", -- $0c768
          51049 => x"00", -- $0c769
          51050 => x"00", -- $0c76a
          51051 => x"00", -- $0c76b
          51052 => x"00", -- $0c76c
          51053 => x"00", -- $0c76d
          51054 => x"00", -- $0c76e
          51055 => x"00", -- $0c76f
          51056 => x"00", -- $0c770
          51057 => x"00", -- $0c771
          51058 => x"00", -- $0c772
          51059 => x"00", -- $0c773
          51060 => x"00", -- $0c774
          51061 => x"00", -- $0c775
          51062 => x"00", -- $0c776
          51063 => x"00", -- $0c777
          51064 => x"00", -- $0c778
          51065 => x"00", -- $0c779
          51066 => x"00", -- $0c77a
          51067 => x"00", -- $0c77b
          51068 => x"00", -- $0c77c
          51069 => x"00", -- $0c77d
          51070 => x"00", -- $0c77e
          51071 => x"00", -- $0c77f
          51072 => x"00", -- $0c780
          51073 => x"00", -- $0c781
          51074 => x"00", -- $0c782
          51075 => x"00", -- $0c783
          51076 => x"00", -- $0c784
          51077 => x"00", -- $0c785
          51078 => x"00", -- $0c786
          51079 => x"00", -- $0c787
          51080 => x"00", -- $0c788
          51081 => x"00", -- $0c789
          51082 => x"00", -- $0c78a
          51083 => x"00", -- $0c78b
          51084 => x"00", -- $0c78c
          51085 => x"00", -- $0c78d
          51086 => x"00", -- $0c78e
          51087 => x"00", -- $0c78f
          51088 => x"00", -- $0c790
          51089 => x"00", -- $0c791
          51090 => x"00", -- $0c792
          51091 => x"00", -- $0c793
          51092 => x"00", -- $0c794
          51093 => x"00", -- $0c795
          51094 => x"00", -- $0c796
          51095 => x"00", -- $0c797
          51096 => x"00", -- $0c798
          51097 => x"00", -- $0c799
          51098 => x"00", -- $0c79a
          51099 => x"00", -- $0c79b
          51100 => x"00", -- $0c79c
          51101 => x"00", -- $0c79d
          51102 => x"00", -- $0c79e
          51103 => x"00", -- $0c79f
          51104 => x"00", -- $0c7a0
          51105 => x"00", -- $0c7a1
          51106 => x"00", -- $0c7a2
          51107 => x"00", -- $0c7a3
          51108 => x"00", -- $0c7a4
          51109 => x"00", -- $0c7a5
          51110 => x"00", -- $0c7a6
          51111 => x"00", -- $0c7a7
          51112 => x"00", -- $0c7a8
          51113 => x"00", -- $0c7a9
          51114 => x"00", -- $0c7aa
          51115 => x"00", -- $0c7ab
          51116 => x"00", -- $0c7ac
          51117 => x"00", -- $0c7ad
          51118 => x"00", -- $0c7ae
          51119 => x"00", -- $0c7af
          51120 => x"00", -- $0c7b0
          51121 => x"00", -- $0c7b1
          51122 => x"00", -- $0c7b2
          51123 => x"00", -- $0c7b3
          51124 => x"00", -- $0c7b4
          51125 => x"00", -- $0c7b5
          51126 => x"00", -- $0c7b6
          51127 => x"00", -- $0c7b7
          51128 => x"00", -- $0c7b8
          51129 => x"00", -- $0c7b9
          51130 => x"00", -- $0c7ba
          51131 => x"00", -- $0c7bb
          51132 => x"00", -- $0c7bc
          51133 => x"00", -- $0c7bd
          51134 => x"00", -- $0c7be
          51135 => x"00", -- $0c7bf
          51136 => x"00", -- $0c7c0
          51137 => x"00", -- $0c7c1
          51138 => x"00", -- $0c7c2
          51139 => x"00", -- $0c7c3
          51140 => x"00", -- $0c7c4
          51141 => x"00", -- $0c7c5
          51142 => x"00", -- $0c7c6
          51143 => x"00", -- $0c7c7
          51144 => x"00", -- $0c7c8
          51145 => x"00", -- $0c7c9
          51146 => x"00", -- $0c7ca
          51147 => x"00", -- $0c7cb
          51148 => x"00", -- $0c7cc
          51149 => x"00", -- $0c7cd
          51150 => x"00", -- $0c7ce
          51151 => x"00", -- $0c7cf
          51152 => x"00", -- $0c7d0
          51153 => x"00", -- $0c7d1
          51154 => x"00", -- $0c7d2
          51155 => x"00", -- $0c7d3
          51156 => x"00", -- $0c7d4
          51157 => x"00", -- $0c7d5
          51158 => x"00", -- $0c7d6
          51159 => x"00", -- $0c7d7
          51160 => x"00", -- $0c7d8
          51161 => x"00", -- $0c7d9
          51162 => x"00", -- $0c7da
          51163 => x"00", -- $0c7db
          51164 => x"00", -- $0c7dc
          51165 => x"00", -- $0c7dd
          51166 => x"00", -- $0c7de
          51167 => x"00", -- $0c7df
          51168 => x"00", -- $0c7e0
          51169 => x"00", -- $0c7e1
          51170 => x"00", -- $0c7e2
          51171 => x"00", -- $0c7e3
          51172 => x"00", -- $0c7e4
          51173 => x"00", -- $0c7e5
          51174 => x"00", -- $0c7e6
          51175 => x"00", -- $0c7e7
          51176 => x"00", -- $0c7e8
          51177 => x"00", -- $0c7e9
          51178 => x"00", -- $0c7ea
          51179 => x"00", -- $0c7eb
          51180 => x"00", -- $0c7ec
          51181 => x"00", -- $0c7ed
          51182 => x"00", -- $0c7ee
          51183 => x"00", -- $0c7ef
          51184 => x"00", -- $0c7f0
          51185 => x"00", -- $0c7f1
          51186 => x"00", -- $0c7f2
          51187 => x"00", -- $0c7f3
          51188 => x"00", -- $0c7f4
          51189 => x"00", -- $0c7f5
          51190 => x"00", -- $0c7f6
          51191 => x"00", -- $0c7f7
          51192 => x"00", -- $0c7f8
          51193 => x"00", -- $0c7f9
          51194 => x"00", -- $0c7fa
          51195 => x"00", -- $0c7fb
          51196 => x"00", -- $0c7fc
          51197 => x"00", -- $0c7fd
          51198 => x"00", -- $0c7fe
          51199 => x"00", -- $0c7ff
          51200 => x"00", -- $0c800
          51201 => x"00", -- $0c801
          51202 => x"00", -- $0c802
          51203 => x"00", -- $0c803
          51204 => x"00", -- $0c804
          51205 => x"00", -- $0c805
          51206 => x"00", -- $0c806
          51207 => x"00", -- $0c807
          51208 => x"00", -- $0c808
          51209 => x"00", -- $0c809
          51210 => x"00", -- $0c80a
          51211 => x"00", -- $0c80b
          51212 => x"00", -- $0c80c
          51213 => x"00", -- $0c80d
          51214 => x"00", -- $0c80e
          51215 => x"00", -- $0c80f
          51216 => x"00", -- $0c810
          51217 => x"00", -- $0c811
          51218 => x"00", -- $0c812
          51219 => x"00", -- $0c813
          51220 => x"00", -- $0c814
          51221 => x"00", -- $0c815
          51222 => x"00", -- $0c816
          51223 => x"00", -- $0c817
          51224 => x"00", -- $0c818
          51225 => x"00", -- $0c819
          51226 => x"00", -- $0c81a
          51227 => x"00", -- $0c81b
          51228 => x"00", -- $0c81c
          51229 => x"00", -- $0c81d
          51230 => x"00", -- $0c81e
          51231 => x"00", -- $0c81f
          51232 => x"00", -- $0c820
          51233 => x"00", -- $0c821
          51234 => x"00", -- $0c822
          51235 => x"00", -- $0c823
          51236 => x"00", -- $0c824
          51237 => x"00", -- $0c825
          51238 => x"00", -- $0c826
          51239 => x"00", -- $0c827
          51240 => x"00", -- $0c828
          51241 => x"00", -- $0c829
          51242 => x"00", -- $0c82a
          51243 => x"00", -- $0c82b
          51244 => x"00", -- $0c82c
          51245 => x"00", -- $0c82d
          51246 => x"00", -- $0c82e
          51247 => x"00", -- $0c82f
          51248 => x"00", -- $0c830
          51249 => x"00", -- $0c831
          51250 => x"00", -- $0c832
          51251 => x"00", -- $0c833
          51252 => x"00", -- $0c834
          51253 => x"00", -- $0c835
          51254 => x"00", -- $0c836
          51255 => x"00", -- $0c837
          51256 => x"00", -- $0c838
          51257 => x"00", -- $0c839
          51258 => x"00", -- $0c83a
          51259 => x"00", -- $0c83b
          51260 => x"00", -- $0c83c
          51261 => x"00", -- $0c83d
          51262 => x"00", -- $0c83e
          51263 => x"00", -- $0c83f
          51264 => x"00", -- $0c840
          51265 => x"00", -- $0c841
          51266 => x"00", -- $0c842
          51267 => x"00", -- $0c843
          51268 => x"00", -- $0c844
          51269 => x"00", -- $0c845
          51270 => x"00", -- $0c846
          51271 => x"00", -- $0c847
          51272 => x"00", -- $0c848
          51273 => x"00", -- $0c849
          51274 => x"00", -- $0c84a
          51275 => x"00", -- $0c84b
          51276 => x"00", -- $0c84c
          51277 => x"00", -- $0c84d
          51278 => x"00", -- $0c84e
          51279 => x"00", -- $0c84f
          51280 => x"00", -- $0c850
          51281 => x"00", -- $0c851
          51282 => x"00", -- $0c852
          51283 => x"00", -- $0c853
          51284 => x"00", -- $0c854
          51285 => x"00", -- $0c855
          51286 => x"00", -- $0c856
          51287 => x"00", -- $0c857
          51288 => x"00", -- $0c858
          51289 => x"00", -- $0c859
          51290 => x"00", -- $0c85a
          51291 => x"00", -- $0c85b
          51292 => x"00", -- $0c85c
          51293 => x"00", -- $0c85d
          51294 => x"00", -- $0c85e
          51295 => x"00", -- $0c85f
          51296 => x"00", -- $0c860
          51297 => x"00", -- $0c861
          51298 => x"00", -- $0c862
          51299 => x"00", -- $0c863
          51300 => x"00", -- $0c864
          51301 => x"00", -- $0c865
          51302 => x"00", -- $0c866
          51303 => x"00", -- $0c867
          51304 => x"00", -- $0c868
          51305 => x"00", -- $0c869
          51306 => x"00", -- $0c86a
          51307 => x"00", -- $0c86b
          51308 => x"00", -- $0c86c
          51309 => x"00", -- $0c86d
          51310 => x"00", -- $0c86e
          51311 => x"00", -- $0c86f
          51312 => x"00", -- $0c870
          51313 => x"00", -- $0c871
          51314 => x"00", -- $0c872
          51315 => x"00", -- $0c873
          51316 => x"00", -- $0c874
          51317 => x"00", -- $0c875
          51318 => x"00", -- $0c876
          51319 => x"00", -- $0c877
          51320 => x"00", -- $0c878
          51321 => x"00", -- $0c879
          51322 => x"00", -- $0c87a
          51323 => x"00", -- $0c87b
          51324 => x"00", -- $0c87c
          51325 => x"00", -- $0c87d
          51326 => x"00", -- $0c87e
          51327 => x"00", -- $0c87f
          51328 => x"00", -- $0c880
          51329 => x"00", -- $0c881
          51330 => x"00", -- $0c882
          51331 => x"00", -- $0c883
          51332 => x"00", -- $0c884
          51333 => x"00", -- $0c885
          51334 => x"00", -- $0c886
          51335 => x"00", -- $0c887
          51336 => x"00", -- $0c888
          51337 => x"00", -- $0c889
          51338 => x"00", -- $0c88a
          51339 => x"00", -- $0c88b
          51340 => x"00", -- $0c88c
          51341 => x"00", -- $0c88d
          51342 => x"00", -- $0c88e
          51343 => x"00", -- $0c88f
          51344 => x"00", -- $0c890
          51345 => x"00", -- $0c891
          51346 => x"00", -- $0c892
          51347 => x"00", -- $0c893
          51348 => x"00", -- $0c894
          51349 => x"00", -- $0c895
          51350 => x"00", -- $0c896
          51351 => x"00", -- $0c897
          51352 => x"00", -- $0c898
          51353 => x"00", -- $0c899
          51354 => x"00", -- $0c89a
          51355 => x"00", -- $0c89b
          51356 => x"00", -- $0c89c
          51357 => x"00", -- $0c89d
          51358 => x"00", -- $0c89e
          51359 => x"00", -- $0c89f
          51360 => x"00", -- $0c8a0
          51361 => x"00", -- $0c8a1
          51362 => x"00", -- $0c8a2
          51363 => x"00", -- $0c8a3
          51364 => x"00", -- $0c8a4
          51365 => x"00", -- $0c8a5
          51366 => x"00", -- $0c8a6
          51367 => x"00", -- $0c8a7
          51368 => x"00", -- $0c8a8
          51369 => x"00", -- $0c8a9
          51370 => x"00", -- $0c8aa
          51371 => x"00", -- $0c8ab
          51372 => x"00", -- $0c8ac
          51373 => x"00", -- $0c8ad
          51374 => x"00", -- $0c8ae
          51375 => x"00", -- $0c8af
          51376 => x"00", -- $0c8b0
          51377 => x"00", -- $0c8b1
          51378 => x"00", -- $0c8b2
          51379 => x"00", -- $0c8b3
          51380 => x"00", -- $0c8b4
          51381 => x"00", -- $0c8b5
          51382 => x"00", -- $0c8b6
          51383 => x"00", -- $0c8b7
          51384 => x"00", -- $0c8b8
          51385 => x"00", -- $0c8b9
          51386 => x"00", -- $0c8ba
          51387 => x"00", -- $0c8bb
          51388 => x"00", -- $0c8bc
          51389 => x"00", -- $0c8bd
          51390 => x"00", -- $0c8be
          51391 => x"00", -- $0c8bf
          51392 => x"00", -- $0c8c0
          51393 => x"00", -- $0c8c1
          51394 => x"00", -- $0c8c2
          51395 => x"00", -- $0c8c3
          51396 => x"00", -- $0c8c4
          51397 => x"00", -- $0c8c5
          51398 => x"00", -- $0c8c6
          51399 => x"00", -- $0c8c7
          51400 => x"00", -- $0c8c8
          51401 => x"00", -- $0c8c9
          51402 => x"00", -- $0c8ca
          51403 => x"00", -- $0c8cb
          51404 => x"00", -- $0c8cc
          51405 => x"00", -- $0c8cd
          51406 => x"00", -- $0c8ce
          51407 => x"00", -- $0c8cf
          51408 => x"00", -- $0c8d0
          51409 => x"00", -- $0c8d1
          51410 => x"00", -- $0c8d2
          51411 => x"00", -- $0c8d3
          51412 => x"00", -- $0c8d4
          51413 => x"00", -- $0c8d5
          51414 => x"00", -- $0c8d6
          51415 => x"00", -- $0c8d7
          51416 => x"00", -- $0c8d8
          51417 => x"00", -- $0c8d9
          51418 => x"00", -- $0c8da
          51419 => x"00", -- $0c8db
          51420 => x"00", -- $0c8dc
          51421 => x"00", -- $0c8dd
          51422 => x"00", -- $0c8de
          51423 => x"00", -- $0c8df
          51424 => x"00", -- $0c8e0
          51425 => x"00", -- $0c8e1
          51426 => x"00", -- $0c8e2
          51427 => x"00", -- $0c8e3
          51428 => x"00", -- $0c8e4
          51429 => x"00", -- $0c8e5
          51430 => x"00", -- $0c8e6
          51431 => x"00", -- $0c8e7
          51432 => x"00", -- $0c8e8
          51433 => x"00", -- $0c8e9
          51434 => x"00", -- $0c8ea
          51435 => x"00", -- $0c8eb
          51436 => x"00", -- $0c8ec
          51437 => x"00", -- $0c8ed
          51438 => x"00", -- $0c8ee
          51439 => x"00", -- $0c8ef
          51440 => x"00", -- $0c8f0
          51441 => x"00", -- $0c8f1
          51442 => x"00", -- $0c8f2
          51443 => x"00", -- $0c8f3
          51444 => x"00", -- $0c8f4
          51445 => x"00", -- $0c8f5
          51446 => x"00", -- $0c8f6
          51447 => x"00", -- $0c8f7
          51448 => x"00", -- $0c8f8
          51449 => x"00", -- $0c8f9
          51450 => x"00", -- $0c8fa
          51451 => x"00", -- $0c8fb
          51452 => x"00", -- $0c8fc
          51453 => x"00", -- $0c8fd
          51454 => x"00", -- $0c8fe
          51455 => x"00", -- $0c8ff
          51456 => x"00", -- $0c900
          51457 => x"00", -- $0c901
          51458 => x"00", -- $0c902
          51459 => x"00", -- $0c903
          51460 => x"00", -- $0c904
          51461 => x"00", -- $0c905
          51462 => x"00", -- $0c906
          51463 => x"00", -- $0c907
          51464 => x"00", -- $0c908
          51465 => x"00", -- $0c909
          51466 => x"00", -- $0c90a
          51467 => x"00", -- $0c90b
          51468 => x"00", -- $0c90c
          51469 => x"00", -- $0c90d
          51470 => x"00", -- $0c90e
          51471 => x"00", -- $0c90f
          51472 => x"00", -- $0c910
          51473 => x"00", -- $0c911
          51474 => x"00", -- $0c912
          51475 => x"00", -- $0c913
          51476 => x"00", -- $0c914
          51477 => x"00", -- $0c915
          51478 => x"00", -- $0c916
          51479 => x"00", -- $0c917
          51480 => x"00", -- $0c918
          51481 => x"00", -- $0c919
          51482 => x"00", -- $0c91a
          51483 => x"00", -- $0c91b
          51484 => x"00", -- $0c91c
          51485 => x"00", -- $0c91d
          51486 => x"00", -- $0c91e
          51487 => x"00", -- $0c91f
          51488 => x"00", -- $0c920
          51489 => x"00", -- $0c921
          51490 => x"00", -- $0c922
          51491 => x"00", -- $0c923
          51492 => x"00", -- $0c924
          51493 => x"00", -- $0c925
          51494 => x"00", -- $0c926
          51495 => x"00", -- $0c927
          51496 => x"00", -- $0c928
          51497 => x"00", -- $0c929
          51498 => x"00", -- $0c92a
          51499 => x"00", -- $0c92b
          51500 => x"00", -- $0c92c
          51501 => x"00", -- $0c92d
          51502 => x"00", -- $0c92e
          51503 => x"00", -- $0c92f
          51504 => x"00", -- $0c930
          51505 => x"00", -- $0c931
          51506 => x"00", -- $0c932
          51507 => x"00", -- $0c933
          51508 => x"00", -- $0c934
          51509 => x"00", -- $0c935
          51510 => x"00", -- $0c936
          51511 => x"00", -- $0c937
          51512 => x"00", -- $0c938
          51513 => x"00", -- $0c939
          51514 => x"00", -- $0c93a
          51515 => x"00", -- $0c93b
          51516 => x"00", -- $0c93c
          51517 => x"00", -- $0c93d
          51518 => x"00", -- $0c93e
          51519 => x"00", -- $0c93f
          51520 => x"00", -- $0c940
          51521 => x"00", -- $0c941
          51522 => x"00", -- $0c942
          51523 => x"00", -- $0c943
          51524 => x"00", -- $0c944
          51525 => x"00", -- $0c945
          51526 => x"00", -- $0c946
          51527 => x"00", -- $0c947
          51528 => x"00", -- $0c948
          51529 => x"00", -- $0c949
          51530 => x"00", -- $0c94a
          51531 => x"00", -- $0c94b
          51532 => x"00", -- $0c94c
          51533 => x"00", -- $0c94d
          51534 => x"00", -- $0c94e
          51535 => x"00", -- $0c94f
          51536 => x"00", -- $0c950
          51537 => x"00", -- $0c951
          51538 => x"00", -- $0c952
          51539 => x"00", -- $0c953
          51540 => x"00", -- $0c954
          51541 => x"00", -- $0c955
          51542 => x"00", -- $0c956
          51543 => x"00", -- $0c957
          51544 => x"00", -- $0c958
          51545 => x"00", -- $0c959
          51546 => x"00", -- $0c95a
          51547 => x"00", -- $0c95b
          51548 => x"00", -- $0c95c
          51549 => x"00", -- $0c95d
          51550 => x"00", -- $0c95e
          51551 => x"00", -- $0c95f
          51552 => x"00", -- $0c960
          51553 => x"00", -- $0c961
          51554 => x"00", -- $0c962
          51555 => x"00", -- $0c963
          51556 => x"00", -- $0c964
          51557 => x"00", -- $0c965
          51558 => x"00", -- $0c966
          51559 => x"00", -- $0c967
          51560 => x"00", -- $0c968
          51561 => x"00", -- $0c969
          51562 => x"00", -- $0c96a
          51563 => x"00", -- $0c96b
          51564 => x"00", -- $0c96c
          51565 => x"00", -- $0c96d
          51566 => x"00", -- $0c96e
          51567 => x"00", -- $0c96f
          51568 => x"00", -- $0c970
          51569 => x"00", -- $0c971
          51570 => x"00", -- $0c972
          51571 => x"00", -- $0c973
          51572 => x"00", -- $0c974
          51573 => x"00", -- $0c975
          51574 => x"00", -- $0c976
          51575 => x"00", -- $0c977
          51576 => x"00", -- $0c978
          51577 => x"00", -- $0c979
          51578 => x"00", -- $0c97a
          51579 => x"00", -- $0c97b
          51580 => x"00", -- $0c97c
          51581 => x"00", -- $0c97d
          51582 => x"00", -- $0c97e
          51583 => x"00", -- $0c97f
          51584 => x"00", -- $0c980
          51585 => x"00", -- $0c981
          51586 => x"00", -- $0c982
          51587 => x"00", -- $0c983
          51588 => x"00", -- $0c984
          51589 => x"00", -- $0c985
          51590 => x"00", -- $0c986
          51591 => x"00", -- $0c987
          51592 => x"00", -- $0c988
          51593 => x"00", -- $0c989
          51594 => x"00", -- $0c98a
          51595 => x"00", -- $0c98b
          51596 => x"00", -- $0c98c
          51597 => x"00", -- $0c98d
          51598 => x"00", -- $0c98e
          51599 => x"00", -- $0c98f
          51600 => x"00", -- $0c990
          51601 => x"00", -- $0c991
          51602 => x"00", -- $0c992
          51603 => x"00", -- $0c993
          51604 => x"00", -- $0c994
          51605 => x"00", -- $0c995
          51606 => x"00", -- $0c996
          51607 => x"00", -- $0c997
          51608 => x"00", -- $0c998
          51609 => x"00", -- $0c999
          51610 => x"00", -- $0c99a
          51611 => x"00", -- $0c99b
          51612 => x"00", -- $0c99c
          51613 => x"00", -- $0c99d
          51614 => x"00", -- $0c99e
          51615 => x"00", -- $0c99f
          51616 => x"00", -- $0c9a0
          51617 => x"00", -- $0c9a1
          51618 => x"00", -- $0c9a2
          51619 => x"00", -- $0c9a3
          51620 => x"00", -- $0c9a4
          51621 => x"00", -- $0c9a5
          51622 => x"00", -- $0c9a6
          51623 => x"00", -- $0c9a7
          51624 => x"00", -- $0c9a8
          51625 => x"00", -- $0c9a9
          51626 => x"00", -- $0c9aa
          51627 => x"00", -- $0c9ab
          51628 => x"00", -- $0c9ac
          51629 => x"00", -- $0c9ad
          51630 => x"00", -- $0c9ae
          51631 => x"00", -- $0c9af
          51632 => x"00", -- $0c9b0
          51633 => x"00", -- $0c9b1
          51634 => x"00", -- $0c9b2
          51635 => x"00", -- $0c9b3
          51636 => x"00", -- $0c9b4
          51637 => x"00", -- $0c9b5
          51638 => x"00", -- $0c9b6
          51639 => x"00", -- $0c9b7
          51640 => x"00", -- $0c9b8
          51641 => x"00", -- $0c9b9
          51642 => x"00", -- $0c9ba
          51643 => x"00", -- $0c9bb
          51644 => x"00", -- $0c9bc
          51645 => x"00", -- $0c9bd
          51646 => x"00", -- $0c9be
          51647 => x"00", -- $0c9bf
          51648 => x"00", -- $0c9c0
          51649 => x"00", -- $0c9c1
          51650 => x"00", -- $0c9c2
          51651 => x"00", -- $0c9c3
          51652 => x"00", -- $0c9c4
          51653 => x"00", -- $0c9c5
          51654 => x"00", -- $0c9c6
          51655 => x"00", -- $0c9c7
          51656 => x"00", -- $0c9c8
          51657 => x"00", -- $0c9c9
          51658 => x"00", -- $0c9ca
          51659 => x"00", -- $0c9cb
          51660 => x"00", -- $0c9cc
          51661 => x"00", -- $0c9cd
          51662 => x"00", -- $0c9ce
          51663 => x"00", -- $0c9cf
          51664 => x"00", -- $0c9d0
          51665 => x"00", -- $0c9d1
          51666 => x"00", -- $0c9d2
          51667 => x"00", -- $0c9d3
          51668 => x"00", -- $0c9d4
          51669 => x"00", -- $0c9d5
          51670 => x"00", -- $0c9d6
          51671 => x"00", -- $0c9d7
          51672 => x"00", -- $0c9d8
          51673 => x"00", -- $0c9d9
          51674 => x"00", -- $0c9da
          51675 => x"00", -- $0c9db
          51676 => x"00", -- $0c9dc
          51677 => x"00", -- $0c9dd
          51678 => x"00", -- $0c9de
          51679 => x"00", -- $0c9df
          51680 => x"00", -- $0c9e0
          51681 => x"00", -- $0c9e1
          51682 => x"00", -- $0c9e2
          51683 => x"00", -- $0c9e3
          51684 => x"00", -- $0c9e4
          51685 => x"00", -- $0c9e5
          51686 => x"00", -- $0c9e6
          51687 => x"00", -- $0c9e7
          51688 => x"00", -- $0c9e8
          51689 => x"00", -- $0c9e9
          51690 => x"00", -- $0c9ea
          51691 => x"00", -- $0c9eb
          51692 => x"00", -- $0c9ec
          51693 => x"00", -- $0c9ed
          51694 => x"00", -- $0c9ee
          51695 => x"00", -- $0c9ef
          51696 => x"00", -- $0c9f0
          51697 => x"00", -- $0c9f1
          51698 => x"00", -- $0c9f2
          51699 => x"00", -- $0c9f3
          51700 => x"00", -- $0c9f4
          51701 => x"00", -- $0c9f5
          51702 => x"00", -- $0c9f6
          51703 => x"00", -- $0c9f7
          51704 => x"00", -- $0c9f8
          51705 => x"00", -- $0c9f9
          51706 => x"00", -- $0c9fa
          51707 => x"00", -- $0c9fb
          51708 => x"00", -- $0c9fc
          51709 => x"00", -- $0c9fd
          51710 => x"00", -- $0c9fe
          51711 => x"00", -- $0c9ff
          51712 => x"00", -- $0ca00
          51713 => x"00", -- $0ca01
          51714 => x"00", -- $0ca02
          51715 => x"00", -- $0ca03
          51716 => x"00", -- $0ca04
          51717 => x"00", -- $0ca05
          51718 => x"00", -- $0ca06
          51719 => x"00", -- $0ca07
          51720 => x"00", -- $0ca08
          51721 => x"00", -- $0ca09
          51722 => x"00", -- $0ca0a
          51723 => x"00", -- $0ca0b
          51724 => x"00", -- $0ca0c
          51725 => x"00", -- $0ca0d
          51726 => x"00", -- $0ca0e
          51727 => x"00", -- $0ca0f
          51728 => x"00", -- $0ca10
          51729 => x"00", -- $0ca11
          51730 => x"00", -- $0ca12
          51731 => x"00", -- $0ca13
          51732 => x"00", -- $0ca14
          51733 => x"00", -- $0ca15
          51734 => x"00", -- $0ca16
          51735 => x"00", -- $0ca17
          51736 => x"00", -- $0ca18
          51737 => x"00", -- $0ca19
          51738 => x"00", -- $0ca1a
          51739 => x"00", -- $0ca1b
          51740 => x"00", -- $0ca1c
          51741 => x"00", -- $0ca1d
          51742 => x"00", -- $0ca1e
          51743 => x"00", -- $0ca1f
          51744 => x"00", -- $0ca20
          51745 => x"00", -- $0ca21
          51746 => x"00", -- $0ca22
          51747 => x"00", -- $0ca23
          51748 => x"00", -- $0ca24
          51749 => x"00", -- $0ca25
          51750 => x"00", -- $0ca26
          51751 => x"00", -- $0ca27
          51752 => x"00", -- $0ca28
          51753 => x"00", -- $0ca29
          51754 => x"00", -- $0ca2a
          51755 => x"00", -- $0ca2b
          51756 => x"00", -- $0ca2c
          51757 => x"00", -- $0ca2d
          51758 => x"00", -- $0ca2e
          51759 => x"00", -- $0ca2f
          51760 => x"00", -- $0ca30
          51761 => x"00", -- $0ca31
          51762 => x"00", -- $0ca32
          51763 => x"00", -- $0ca33
          51764 => x"00", -- $0ca34
          51765 => x"00", -- $0ca35
          51766 => x"00", -- $0ca36
          51767 => x"00", -- $0ca37
          51768 => x"00", -- $0ca38
          51769 => x"00", -- $0ca39
          51770 => x"00", -- $0ca3a
          51771 => x"00", -- $0ca3b
          51772 => x"00", -- $0ca3c
          51773 => x"00", -- $0ca3d
          51774 => x"00", -- $0ca3e
          51775 => x"00", -- $0ca3f
          51776 => x"00", -- $0ca40
          51777 => x"00", -- $0ca41
          51778 => x"00", -- $0ca42
          51779 => x"00", -- $0ca43
          51780 => x"00", -- $0ca44
          51781 => x"00", -- $0ca45
          51782 => x"00", -- $0ca46
          51783 => x"00", -- $0ca47
          51784 => x"00", -- $0ca48
          51785 => x"00", -- $0ca49
          51786 => x"00", -- $0ca4a
          51787 => x"00", -- $0ca4b
          51788 => x"00", -- $0ca4c
          51789 => x"00", -- $0ca4d
          51790 => x"00", -- $0ca4e
          51791 => x"00", -- $0ca4f
          51792 => x"00", -- $0ca50
          51793 => x"00", -- $0ca51
          51794 => x"00", -- $0ca52
          51795 => x"00", -- $0ca53
          51796 => x"00", -- $0ca54
          51797 => x"00", -- $0ca55
          51798 => x"00", -- $0ca56
          51799 => x"00", -- $0ca57
          51800 => x"00", -- $0ca58
          51801 => x"00", -- $0ca59
          51802 => x"00", -- $0ca5a
          51803 => x"00", -- $0ca5b
          51804 => x"00", -- $0ca5c
          51805 => x"00", -- $0ca5d
          51806 => x"00", -- $0ca5e
          51807 => x"00", -- $0ca5f
          51808 => x"00", -- $0ca60
          51809 => x"00", -- $0ca61
          51810 => x"00", -- $0ca62
          51811 => x"00", -- $0ca63
          51812 => x"00", -- $0ca64
          51813 => x"00", -- $0ca65
          51814 => x"00", -- $0ca66
          51815 => x"00", -- $0ca67
          51816 => x"00", -- $0ca68
          51817 => x"00", -- $0ca69
          51818 => x"00", -- $0ca6a
          51819 => x"00", -- $0ca6b
          51820 => x"00", -- $0ca6c
          51821 => x"00", -- $0ca6d
          51822 => x"00", -- $0ca6e
          51823 => x"00", -- $0ca6f
          51824 => x"00", -- $0ca70
          51825 => x"00", -- $0ca71
          51826 => x"00", -- $0ca72
          51827 => x"00", -- $0ca73
          51828 => x"00", -- $0ca74
          51829 => x"00", -- $0ca75
          51830 => x"00", -- $0ca76
          51831 => x"00", -- $0ca77
          51832 => x"00", -- $0ca78
          51833 => x"00", -- $0ca79
          51834 => x"00", -- $0ca7a
          51835 => x"00", -- $0ca7b
          51836 => x"00", -- $0ca7c
          51837 => x"00", -- $0ca7d
          51838 => x"00", -- $0ca7e
          51839 => x"00", -- $0ca7f
          51840 => x"00", -- $0ca80
          51841 => x"00", -- $0ca81
          51842 => x"00", -- $0ca82
          51843 => x"00", -- $0ca83
          51844 => x"00", -- $0ca84
          51845 => x"00", -- $0ca85
          51846 => x"00", -- $0ca86
          51847 => x"00", -- $0ca87
          51848 => x"00", -- $0ca88
          51849 => x"00", -- $0ca89
          51850 => x"00", -- $0ca8a
          51851 => x"00", -- $0ca8b
          51852 => x"00", -- $0ca8c
          51853 => x"00", -- $0ca8d
          51854 => x"00", -- $0ca8e
          51855 => x"00", -- $0ca8f
          51856 => x"00", -- $0ca90
          51857 => x"00", -- $0ca91
          51858 => x"00", -- $0ca92
          51859 => x"00", -- $0ca93
          51860 => x"00", -- $0ca94
          51861 => x"00", -- $0ca95
          51862 => x"00", -- $0ca96
          51863 => x"00", -- $0ca97
          51864 => x"00", -- $0ca98
          51865 => x"00", -- $0ca99
          51866 => x"00", -- $0ca9a
          51867 => x"00", -- $0ca9b
          51868 => x"00", -- $0ca9c
          51869 => x"00", -- $0ca9d
          51870 => x"00", -- $0ca9e
          51871 => x"00", -- $0ca9f
          51872 => x"00", -- $0caa0
          51873 => x"00", -- $0caa1
          51874 => x"00", -- $0caa2
          51875 => x"00", -- $0caa3
          51876 => x"00", -- $0caa4
          51877 => x"00", -- $0caa5
          51878 => x"00", -- $0caa6
          51879 => x"00", -- $0caa7
          51880 => x"00", -- $0caa8
          51881 => x"00", -- $0caa9
          51882 => x"00", -- $0caaa
          51883 => x"00", -- $0caab
          51884 => x"00", -- $0caac
          51885 => x"00", -- $0caad
          51886 => x"00", -- $0caae
          51887 => x"00", -- $0caaf
          51888 => x"00", -- $0cab0
          51889 => x"00", -- $0cab1
          51890 => x"00", -- $0cab2
          51891 => x"00", -- $0cab3
          51892 => x"00", -- $0cab4
          51893 => x"00", -- $0cab5
          51894 => x"00", -- $0cab6
          51895 => x"00", -- $0cab7
          51896 => x"00", -- $0cab8
          51897 => x"00", -- $0cab9
          51898 => x"00", -- $0caba
          51899 => x"00", -- $0cabb
          51900 => x"00", -- $0cabc
          51901 => x"00", -- $0cabd
          51902 => x"00", -- $0cabe
          51903 => x"00", -- $0cabf
          51904 => x"00", -- $0cac0
          51905 => x"00", -- $0cac1
          51906 => x"00", -- $0cac2
          51907 => x"00", -- $0cac3
          51908 => x"00", -- $0cac4
          51909 => x"00", -- $0cac5
          51910 => x"00", -- $0cac6
          51911 => x"00", -- $0cac7
          51912 => x"00", -- $0cac8
          51913 => x"00", -- $0cac9
          51914 => x"00", -- $0caca
          51915 => x"00", -- $0cacb
          51916 => x"00", -- $0cacc
          51917 => x"00", -- $0cacd
          51918 => x"00", -- $0cace
          51919 => x"00", -- $0cacf
          51920 => x"00", -- $0cad0
          51921 => x"00", -- $0cad1
          51922 => x"00", -- $0cad2
          51923 => x"00", -- $0cad3
          51924 => x"00", -- $0cad4
          51925 => x"00", -- $0cad5
          51926 => x"00", -- $0cad6
          51927 => x"00", -- $0cad7
          51928 => x"00", -- $0cad8
          51929 => x"00", -- $0cad9
          51930 => x"00", -- $0cada
          51931 => x"00", -- $0cadb
          51932 => x"00", -- $0cadc
          51933 => x"00", -- $0cadd
          51934 => x"00", -- $0cade
          51935 => x"00", -- $0cadf
          51936 => x"00", -- $0cae0
          51937 => x"00", -- $0cae1
          51938 => x"00", -- $0cae2
          51939 => x"00", -- $0cae3
          51940 => x"00", -- $0cae4
          51941 => x"00", -- $0cae5
          51942 => x"00", -- $0cae6
          51943 => x"00", -- $0cae7
          51944 => x"00", -- $0cae8
          51945 => x"00", -- $0cae9
          51946 => x"00", -- $0caea
          51947 => x"00", -- $0caeb
          51948 => x"00", -- $0caec
          51949 => x"00", -- $0caed
          51950 => x"00", -- $0caee
          51951 => x"00", -- $0caef
          51952 => x"00", -- $0caf0
          51953 => x"00", -- $0caf1
          51954 => x"00", -- $0caf2
          51955 => x"00", -- $0caf3
          51956 => x"00", -- $0caf4
          51957 => x"00", -- $0caf5
          51958 => x"00", -- $0caf6
          51959 => x"00", -- $0caf7
          51960 => x"00", -- $0caf8
          51961 => x"00", -- $0caf9
          51962 => x"00", -- $0cafa
          51963 => x"00", -- $0cafb
          51964 => x"00", -- $0cafc
          51965 => x"00", -- $0cafd
          51966 => x"00", -- $0cafe
          51967 => x"00", -- $0caff
          51968 => x"00", -- $0cb00
          51969 => x"00", -- $0cb01
          51970 => x"00", -- $0cb02
          51971 => x"00", -- $0cb03
          51972 => x"00", -- $0cb04
          51973 => x"00", -- $0cb05
          51974 => x"00", -- $0cb06
          51975 => x"00", -- $0cb07
          51976 => x"00", -- $0cb08
          51977 => x"00", -- $0cb09
          51978 => x"00", -- $0cb0a
          51979 => x"00", -- $0cb0b
          51980 => x"00", -- $0cb0c
          51981 => x"00", -- $0cb0d
          51982 => x"00", -- $0cb0e
          51983 => x"00", -- $0cb0f
          51984 => x"00", -- $0cb10
          51985 => x"00", -- $0cb11
          51986 => x"00", -- $0cb12
          51987 => x"00", -- $0cb13
          51988 => x"00", -- $0cb14
          51989 => x"00", -- $0cb15
          51990 => x"00", -- $0cb16
          51991 => x"00", -- $0cb17
          51992 => x"00", -- $0cb18
          51993 => x"00", -- $0cb19
          51994 => x"00", -- $0cb1a
          51995 => x"00", -- $0cb1b
          51996 => x"00", -- $0cb1c
          51997 => x"00", -- $0cb1d
          51998 => x"00", -- $0cb1e
          51999 => x"00", -- $0cb1f
          52000 => x"00", -- $0cb20
          52001 => x"00", -- $0cb21
          52002 => x"00", -- $0cb22
          52003 => x"00", -- $0cb23
          52004 => x"00", -- $0cb24
          52005 => x"00", -- $0cb25
          52006 => x"00", -- $0cb26
          52007 => x"00", -- $0cb27
          52008 => x"00", -- $0cb28
          52009 => x"00", -- $0cb29
          52010 => x"00", -- $0cb2a
          52011 => x"00", -- $0cb2b
          52012 => x"00", -- $0cb2c
          52013 => x"00", -- $0cb2d
          52014 => x"00", -- $0cb2e
          52015 => x"00", -- $0cb2f
          52016 => x"00", -- $0cb30
          52017 => x"00", -- $0cb31
          52018 => x"00", -- $0cb32
          52019 => x"00", -- $0cb33
          52020 => x"00", -- $0cb34
          52021 => x"00", -- $0cb35
          52022 => x"00", -- $0cb36
          52023 => x"00", -- $0cb37
          52024 => x"00", -- $0cb38
          52025 => x"00", -- $0cb39
          52026 => x"00", -- $0cb3a
          52027 => x"00", -- $0cb3b
          52028 => x"00", -- $0cb3c
          52029 => x"00", -- $0cb3d
          52030 => x"00", -- $0cb3e
          52031 => x"00", -- $0cb3f
          52032 => x"00", -- $0cb40
          52033 => x"00", -- $0cb41
          52034 => x"00", -- $0cb42
          52035 => x"00", -- $0cb43
          52036 => x"00", -- $0cb44
          52037 => x"00", -- $0cb45
          52038 => x"00", -- $0cb46
          52039 => x"00", -- $0cb47
          52040 => x"00", -- $0cb48
          52041 => x"00", -- $0cb49
          52042 => x"00", -- $0cb4a
          52043 => x"00", -- $0cb4b
          52044 => x"00", -- $0cb4c
          52045 => x"00", -- $0cb4d
          52046 => x"00", -- $0cb4e
          52047 => x"00", -- $0cb4f
          52048 => x"00", -- $0cb50
          52049 => x"00", -- $0cb51
          52050 => x"00", -- $0cb52
          52051 => x"00", -- $0cb53
          52052 => x"00", -- $0cb54
          52053 => x"00", -- $0cb55
          52054 => x"00", -- $0cb56
          52055 => x"00", -- $0cb57
          52056 => x"00", -- $0cb58
          52057 => x"00", -- $0cb59
          52058 => x"00", -- $0cb5a
          52059 => x"00", -- $0cb5b
          52060 => x"00", -- $0cb5c
          52061 => x"00", -- $0cb5d
          52062 => x"00", -- $0cb5e
          52063 => x"00", -- $0cb5f
          52064 => x"00", -- $0cb60
          52065 => x"00", -- $0cb61
          52066 => x"00", -- $0cb62
          52067 => x"00", -- $0cb63
          52068 => x"00", -- $0cb64
          52069 => x"00", -- $0cb65
          52070 => x"00", -- $0cb66
          52071 => x"00", -- $0cb67
          52072 => x"00", -- $0cb68
          52073 => x"00", -- $0cb69
          52074 => x"00", -- $0cb6a
          52075 => x"00", -- $0cb6b
          52076 => x"00", -- $0cb6c
          52077 => x"00", -- $0cb6d
          52078 => x"00", -- $0cb6e
          52079 => x"00", -- $0cb6f
          52080 => x"00", -- $0cb70
          52081 => x"00", -- $0cb71
          52082 => x"00", -- $0cb72
          52083 => x"00", -- $0cb73
          52084 => x"00", -- $0cb74
          52085 => x"00", -- $0cb75
          52086 => x"00", -- $0cb76
          52087 => x"00", -- $0cb77
          52088 => x"00", -- $0cb78
          52089 => x"00", -- $0cb79
          52090 => x"00", -- $0cb7a
          52091 => x"00", -- $0cb7b
          52092 => x"00", -- $0cb7c
          52093 => x"00", -- $0cb7d
          52094 => x"00", -- $0cb7e
          52095 => x"00", -- $0cb7f
          52096 => x"00", -- $0cb80
          52097 => x"00", -- $0cb81
          52098 => x"00", -- $0cb82
          52099 => x"00", -- $0cb83
          52100 => x"00", -- $0cb84
          52101 => x"00", -- $0cb85
          52102 => x"00", -- $0cb86
          52103 => x"00", -- $0cb87
          52104 => x"00", -- $0cb88
          52105 => x"00", -- $0cb89
          52106 => x"00", -- $0cb8a
          52107 => x"00", -- $0cb8b
          52108 => x"00", -- $0cb8c
          52109 => x"00", -- $0cb8d
          52110 => x"00", -- $0cb8e
          52111 => x"00", -- $0cb8f
          52112 => x"00", -- $0cb90
          52113 => x"00", -- $0cb91
          52114 => x"00", -- $0cb92
          52115 => x"00", -- $0cb93
          52116 => x"00", -- $0cb94
          52117 => x"00", -- $0cb95
          52118 => x"00", -- $0cb96
          52119 => x"00", -- $0cb97
          52120 => x"00", -- $0cb98
          52121 => x"00", -- $0cb99
          52122 => x"00", -- $0cb9a
          52123 => x"00", -- $0cb9b
          52124 => x"00", -- $0cb9c
          52125 => x"00", -- $0cb9d
          52126 => x"00", -- $0cb9e
          52127 => x"00", -- $0cb9f
          52128 => x"00", -- $0cba0
          52129 => x"00", -- $0cba1
          52130 => x"00", -- $0cba2
          52131 => x"00", -- $0cba3
          52132 => x"00", -- $0cba4
          52133 => x"00", -- $0cba5
          52134 => x"00", -- $0cba6
          52135 => x"00", -- $0cba7
          52136 => x"00", -- $0cba8
          52137 => x"00", -- $0cba9
          52138 => x"00", -- $0cbaa
          52139 => x"00", -- $0cbab
          52140 => x"00", -- $0cbac
          52141 => x"00", -- $0cbad
          52142 => x"00", -- $0cbae
          52143 => x"00", -- $0cbaf
          52144 => x"00", -- $0cbb0
          52145 => x"00", -- $0cbb1
          52146 => x"00", -- $0cbb2
          52147 => x"00", -- $0cbb3
          52148 => x"00", -- $0cbb4
          52149 => x"00", -- $0cbb5
          52150 => x"00", -- $0cbb6
          52151 => x"00", -- $0cbb7
          52152 => x"00", -- $0cbb8
          52153 => x"00", -- $0cbb9
          52154 => x"00", -- $0cbba
          52155 => x"00", -- $0cbbb
          52156 => x"00", -- $0cbbc
          52157 => x"00", -- $0cbbd
          52158 => x"00", -- $0cbbe
          52159 => x"00", -- $0cbbf
          52160 => x"00", -- $0cbc0
          52161 => x"00", -- $0cbc1
          52162 => x"00", -- $0cbc2
          52163 => x"00", -- $0cbc3
          52164 => x"00", -- $0cbc4
          52165 => x"00", -- $0cbc5
          52166 => x"00", -- $0cbc6
          52167 => x"00", -- $0cbc7
          52168 => x"00", -- $0cbc8
          52169 => x"00", -- $0cbc9
          52170 => x"00", -- $0cbca
          52171 => x"00", -- $0cbcb
          52172 => x"00", -- $0cbcc
          52173 => x"00", -- $0cbcd
          52174 => x"00", -- $0cbce
          52175 => x"00", -- $0cbcf
          52176 => x"00", -- $0cbd0
          52177 => x"00", -- $0cbd1
          52178 => x"00", -- $0cbd2
          52179 => x"00", -- $0cbd3
          52180 => x"00", -- $0cbd4
          52181 => x"00", -- $0cbd5
          52182 => x"00", -- $0cbd6
          52183 => x"00", -- $0cbd7
          52184 => x"00", -- $0cbd8
          52185 => x"00", -- $0cbd9
          52186 => x"00", -- $0cbda
          52187 => x"00", -- $0cbdb
          52188 => x"00", -- $0cbdc
          52189 => x"00", -- $0cbdd
          52190 => x"00", -- $0cbde
          52191 => x"00", -- $0cbdf
          52192 => x"00", -- $0cbe0
          52193 => x"00", -- $0cbe1
          52194 => x"00", -- $0cbe2
          52195 => x"00", -- $0cbe3
          52196 => x"00", -- $0cbe4
          52197 => x"00", -- $0cbe5
          52198 => x"00", -- $0cbe6
          52199 => x"00", -- $0cbe7
          52200 => x"00", -- $0cbe8
          52201 => x"00", -- $0cbe9
          52202 => x"00", -- $0cbea
          52203 => x"00", -- $0cbeb
          52204 => x"00", -- $0cbec
          52205 => x"00", -- $0cbed
          52206 => x"00", -- $0cbee
          52207 => x"00", -- $0cbef
          52208 => x"00", -- $0cbf0
          52209 => x"00", -- $0cbf1
          52210 => x"00", -- $0cbf2
          52211 => x"00", -- $0cbf3
          52212 => x"00", -- $0cbf4
          52213 => x"00", -- $0cbf5
          52214 => x"00", -- $0cbf6
          52215 => x"00", -- $0cbf7
          52216 => x"00", -- $0cbf8
          52217 => x"00", -- $0cbf9
          52218 => x"00", -- $0cbfa
          52219 => x"00", -- $0cbfb
          52220 => x"00", -- $0cbfc
          52221 => x"00", -- $0cbfd
          52222 => x"00", -- $0cbfe
          52223 => x"00", -- $0cbff
          52224 => x"00", -- $0cc00
          52225 => x"00", -- $0cc01
          52226 => x"00", -- $0cc02
          52227 => x"00", -- $0cc03
          52228 => x"00", -- $0cc04
          52229 => x"00", -- $0cc05
          52230 => x"00", -- $0cc06
          52231 => x"00", -- $0cc07
          52232 => x"00", -- $0cc08
          52233 => x"00", -- $0cc09
          52234 => x"00", -- $0cc0a
          52235 => x"00", -- $0cc0b
          52236 => x"00", -- $0cc0c
          52237 => x"00", -- $0cc0d
          52238 => x"00", -- $0cc0e
          52239 => x"00", -- $0cc0f
          52240 => x"00", -- $0cc10
          52241 => x"00", -- $0cc11
          52242 => x"00", -- $0cc12
          52243 => x"00", -- $0cc13
          52244 => x"00", -- $0cc14
          52245 => x"00", -- $0cc15
          52246 => x"00", -- $0cc16
          52247 => x"00", -- $0cc17
          52248 => x"00", -- $0cc18
          52249 => x"00", -- $0cc19
          52250 => x"00", -- $0cc1a
          52251 => x"00", -- $0cc1b
          52252 => x"00", -- $0cc1c
          52253 => x"00", -- $0cc1d
          52254 => x"00", -- $0cc1e
          52255 => x"00", -- $0cc1f
          52256 => x"00", -- $0cc20
          52257 => x"00", -- $0cc21
          52258 => x"00", -- $0cc22
          52259 => x"00", -- $0cc23
          52260 => x"00", -- $0cc24
          52261 => x"00", -- $0cc25
          52262 => x"00", -- $0cc26
          52263 => x"00", -- $0cc27
          52264 => x"00", -- $0cc28
          52265 => x"00", -- $0cc29
          52266 => x"00", -- $0cc2a
          52267 => x"00", -- $0cc2b
          52268 => x"00", -- $0cc2c
          52269 => x"00", -- $0cc2d
          52270 => x"00", -- $0cc2e
          52271 => x"00", -- $0cc2f
          52272 => x"00", -- $0cc30
          52273 => x"00", -- $0cc31
          52274 => x"00", -- $0cc32
          52275 => x"00", -- $0cc33
          52276 => x"00", -- $0cc34
          52277 => x"00", -- $0cc35
          52278 => x"00", -- $0cc36
          52279 => x"00", -- $0cc37
          52280 => x"00", -- $0cc38
          52281 => x"00", -- $0cc39
          52282 => x"00", -- $0cc3a
          52283 => x"00", -- $0cc3b
          52284 => x"00", -- $0cc3c
          52285 => x"00", -- $0cc3d
          52286 => x"00", -- $0cc3e
          52287 => x"00", -- $0cc3f
          52288 => x"00", -- $0cc40
          52289 => x"00", -- $0cc41
          52290 => x"00", -- $0cc42
          52291 => x"00", -- $0cc43
          52292 => x"00", -- $0cc44
          52293 => x"00", -- $0cc45
          52294 => x"00", -- $0cc46
          52295 => x"00", -- $0cc47
          52296 => x"00", -- $0cc48
          52297 => x"00", -- $0cc49
          52298 => x"00", -- $0cc4a
          52299 => x"00", -- $0cc4b
          52300 => x"00", -- $0cc4c
          52301 => x"00", -- $0cc4d
          52302 => x"00", -- $0cc4e
          52303 => x"00", -- $0cc4f
          52304 => x"00", -- $0cc50
          52305 => x"00", -- $0cc51
          52306 => x"00", -- $0cc52
          52307 => x"00", -- $0cc53
          52308 => x"00", -- $0cc54
          52309 => x"00", -- $0cc55
          52310 => x"00", -- $0cc56
          52311 => x"00", -- $0cc57
          52312 => x"00", -- $0cc58
          52313 => x"00", -- $0cc59
          52314 => x"00", -- $0cc5a
          52315 => x"00", -- $0cc5b
          52316 => x"00", -- $0cc5c
          52317 => x"00", -- $0cc5d
          52318 => x"00", -- $0cc5e
          52319 => x"00", -- $0cc5f
          52320 => x"00", -- $0cc60
          52321 => x"00", -- $0cc61
          52322 => x"00", -- $0cc62
          52323 => x"00", -- $0cc63
          52324 => x"00", -- $0cc64
          52325 => x"00", -- $0cc65
          52326 => x"00", -- $0cc66
          52327 => x"00", -- $0cc67
          52328 => x"00", -- $0cc68
          52329 => x"00", -- $0cc69
          52330 => x"00", -- $0cc6a
          52331 => x"00", -- $0cc6b
          52332 => x"00", -- $0cc6c
          52333 => x"00", -- $0cc6d
          52334 => x"00", -- $0cc6e
          52335 => x"00", -- $0cc6f
          52336 => x"00", -- $0cc70
          52337 => x"00", -- $0cc71
          52338 => x"00", -- $0cc72
          52339 => x"00", -- $0cc73
          52340 => x"00", -- $0cc74
          52341 => x"00", -- $0cc75
          52342 => x"00", -- $0cc76
          52343 => x"00", -- $0cc77
          52344 => x"00", -- $0cc78
          52345 => x"00", -- $0cc79
          52346 => x"00", -- $0cc7a
          52347 => x"00", -- $0cc7b
          52348 => x"00", -- $0cc7c
          52349 => x"00", -- $0cc7d
          52350 => x"00", -- $0cc7e
          52351 => x"00", -- $0cc7f
          52352 => x"00", -- $0cc80
          52353 => x"00", -- $0cc81
          52354 => x"00", -- $0cc82
          52355 => x"00", -- $0cc83
          52356 => x"00", -- $0cc84
          52357 => x"00", -- $0cc85
          52358 => x"00", -- $0cc86
          52359 => x"00", -- $0cc87
          52360 => x"00", -- $0cc88
          52361 => x"00", -- $0cc89
          52362 => x"00", -- $0cc8a
          52363 => x"00", -- $0cc8b
          52364 => x"00", -- $0cc8c
          52365 => x"00", -- $0cc8d
          52366 => x"00", -- $0cc8e
          52367 => x"00", -- $0cc8f
          52368 => x"00", -- $0cc90
          52369 => x"00", -- $0cc91
          52370 => x"00", -- $0cc92
          52371 => x"00", -- $0cc93
          52372 => x"00", -- $0cc94
          52373 => x"00", -- $0cc95
          52374 => x"00", -- $0cc96
          52375 => x"00", -- $0cc97
          52376 => x"00", -- $0cc98
          52377 => x"00", -- $0cc99
          52378 => x"00", -- $0cc9a
          52379 => x"00", -- $0cc9b
          52380 => x"00", -- $0cc9c
          52381 => x"00", -- $0cc9d
          52382 => x"00", -- $0cc9e
          52383 => x"00", -- $0cc9f
          52384 => x"00", -- $0cca0
          52385 => x"00", -- $0cca1
          52386 => x"00", -- $0cca2
          52387 => x"00", -- $0cca3
          52388 => x"00", -- $0cca4
          52389 => x"00", -- $0cca5
          52390 => x"00", -- $0cca6
          52391 => x"00", -- $0cca7
          52392 => x"00", -- $0cca8
          52393 => x"00", -- $0cca9
          52394 => x"00", -- $0ccaa
          52395 => x"00", -- $0ccab
          52396 => x"00", -- $0ccac
          52397 => x"00", -- $0ccad
          52398 => x"00", -- $0ccae
          52399 => x"00", -- $0ccaf
          52400 => x"00", -- $0ccb0
          52401 => x"00", -- $0ccb1
          52402 => x"00", -- $0ccb2
          52403 => x"00", -- $0ccb3
          52404 => x"00", -- $0ccb4
          52405 => x"00", -- $0ccb5
          52406 => x"00", -- $0ccb6
          52407 => x"00", -- $0ccb7
          52408 => x"00", -- $0ccb8
          52409 => x"00", -- $0ccb9
          52410 => x"00", -- $0ccba
          52411 => x"00", -- $0ccbb
          52412 => x"00", -- $0ccbc
          52413 => x"00", -- $0ccbd
          52414 => x"00", -- $0ccbe
          52415 => x"00", -- $0ccbf
          52416 => x"00", -- $0ccc0
          52417 => x"00", -- $0ccc1
          52418 => x"00", -- $0ccc2
          52419 => x"00", -- $0ccc3
          52420 => x"00", -- $0ccc4
          52421 => x"00", -- $0ccc5
          52422 => x"00", -- $0ccc6
          52423 => x"00", -- $0ccc7
          52424 => x"00", -- $0ccc8
          52425 => x"00", -- $0ccc9
          52426 => x"00", -- $0ccca
          52427 => x"00", -- $0cccb
          52428 => x"00", -- $0cccc
          52429 => x"00", -- $0cccd
          52430 => x"00", -- $0ccce
          52431 => x"00", -- $0cccf
          52432 => x"00", -- $0ccd0
          52433 => x"00", -- $0ccd1
          52434 => x"00", -- $0ccd2
          52435 => x"00", -- $0ccd3
          52436 => x"00", -- $0ccd4
          52437 => x"00", -- $0ccd5
          52438 => x"00", -- $0ccd6
          52439 => x"00", -- $0ccd7
          52440 => x"00", -- $0ccd8
          52441 => x"00", -- $0ccd9
          52442 => x"00", -- $0ccda
          52443 => x"00", -- $0ccdb
          52444 => x"00", -- $0ccdc
          52445 => x"00", -- $0ccdd
          52446 => x"00", -- $0ccde
          52447 => x"00", -- $0ccdf
          52448 => x"00", -- $0cce0
          52449 => x"00", -- $0cce1
          52450 => x"00", -- $0cce2
          52451 => x"00", -- $0cce3
          52452 => x"00", -- $0cce4
          52453 => x"00", -- $0cce5
          52454 => x"00", -- $0cce6
          52455 => x"00", -- $0cce7
          52456 => x"00", -- $0cce8
          52457 => x"00", -- $0cce9
          52458 => x"00", -- $0ccea
          52459 => x"00", -- $0cceb
          52460 => x"00", -- $0ccec
          52461 => x"00", -- $0cced
          52462 => x"00", -- $0ccee
          52463 => x"00", -- $0ccef
          52464 => x"00", -- $0ccf0
          52465 => x"00", -- $0ccf1
          52466 => x"00", -- $0ccf2
          52467 => x"00", -- $0ccf3
          52468 => x"00", -- $0ccf4
          52469 => x"00", -- $0ccf5
          52470 => x"00", -- $0ccf6
          52471 => x"00", -- $0ccf7
          52472 => x"00", -- $0ccf8
          52473 => x"00", -- $0ccf9
          52474 => x"00", -- $0ccfa
          52475 => x"00", -- $0ccfb
          52476 => x"00", -- $0ccfc
          52477 => x"00", -- $0ccfd
          52478 => x"00", -- $0ccfe
          52479 => x"00", -- $0ccff
          52480 => x"00", -- $0cd00
          52481 => x"00", -- $0cd01
          52482 => x"00", -- $0cd02
          52483 => x"00", -- $0cd03
          52484 => x"00", -- $0cd04
          52485 => x"00", -- $0cd05
          52486 => x"00", -- $0cd06
          52487 => x"00", -- $0cd07
          52488 => x"00", -- $0cd08
          52489 => x"00", -- $0cd09
          52490 => x"00", -- $0cd0a
          52491 => x"00", -- $0cd0b
          52492 => x"00", -- $0cd0c
          52493 => x"00", -- $0cd0d
          52494 => x"00", -- $0cd0e
          52495 => x"00", -- $0cd0f
          52496 => x"00", -- $0cd10
          52497 => x"00", -- $0cd11
          52498 => x"00", -- $0cd12
          52499 => x"00", -- $0cd13
          52500 => x"00", -- $0cd14
          52501 => x"00", -- $0cd15
          52502 => x"00", -- $0cd16
          52503 => x"00", -- $0cd17
          52504 => x"00", -- $0cd18
          52505 => x"00", -- $0cd19
          52506 => x"00", -- $0cd1a
          52507 => x"00", -- $0cd1b
          52508 => x"00", -- $0cd1c
          52509 => x"00", -- $0cd1d
          52510 => x"00", -- $0cd1e
          52511 => x"00", -- $0cd1f
          52512 => x"00", -- $0cd20
          52513 => x"00", -- $0cd21
          52514 => x"00", -- $0cd22
          52515 => x"00", -- $0cd23
          52516 => x"00", -- $0cd24
          52517 => x"00", -- $0cd25
          52518 => x"00", -- $0cd26
          52519 => x"00", -- $0cd27
          52520 => x"00", -- $0cd28
          52521 => x"00", -- $0cd29
          52522 => x"00", -- $0cd2a
          52523 => x"00", -- $0cd2b
          52524 => x"00", -- $0cd2c
          52525 => x"00", -- $0cd2d
          52526 => x"00", -- $0cd2e
          52527 => x"00", -- $0cd2f
          52528 => x"00", -- $0cd30
          52529 => x"00", -- $0cd31
          52530 => x"00", -- $0cd32
          52531 => x"00", -- $0cd33
          52532 => x"00", -- $0cd34
          52533 => x"00", -- $0cd35
          52534 => x"00", -- $0cd36
          52535 => x"00", -- $0cd37
          52536 => x"00", -- $0cd38
          52537 => x"00", -- $0cd39
          52538 => x"00", -- $0cd3a
          52539 => x"00", -- $0cd3b
          52540 => x"00", -- $0cd3c
          52541 => x"00", -- $0cd3d
          52542 => x"00", -- $0cd3e
          52543 => x"00", -- $0cd3f
          52544 => x"00", -- $0cd40
          52545 => x"00", -- $0cd41
          52546 => x"00", -- $0cd42
          52547 => x"00", -- $0cd43
          52548 => x"00", -- $0cd44
          52549 => x"00", -- $0cd45
          52550 => x"00", -- $0cd46
          52551 => x"00", -- $0cd47
          52552 => x"00", -- $0cd48
          52553 => x"00", -- $0cd49
          52554 => x"00", -- $0cd4a
          52555 => x"00", -- $0cd4b
          52556 => x"00", -- $0cd4c
          52557 => x"00", -- $0cd4d
          52558 => x"00", -- $0cd4e
          52559 => x"00", -- $0cd4f
          52560 => x"00", -- $0cd50
          52561 => x"00", -- $0cd51
          52562 => x"00", -- $0cd52
          52563 => x"00", -- $0cd53
          52564 => x"00", -- $0cd54
          52565 => x"00", -- $0cd55
          52566 => x"00", -- $0cd56
          52567 => x"00", -- $0cd57
          52568 => x"00", -- $0cd58
          52569 => x"00", -- $0cd59
          52570 => x"00", -- $0cd5a
          52571 => x"00", -- $0cd5b
          52572 => x"00", -- $0cd5c
          52573 => x"00", -- $0cd5d
          52574 => x"00", -- $0cd5e
          52575 => x"00", -- $0cd5f
          52576 => x"00", -- $0cd60
          52577 => x"00", -- $0cd61
          52578 => x"00", -- $0cd62
          52579 => x"00", -- $0cd63
          52580 => x"00", -- $0cd64
          52581 => x"00", -- $0cd65
          52582 => x"00", -- $0cd66
          52583 => x"00", -- $0cd67
          52584 => x"00", -- $0cd68
          52585 => x"00", -- $0cd69
          52586 => x"00", -- $0cd6a
          52587 => x"00", -- $0cd6b
          52588 => x"00", -- $0cd6c
          52589 => x"00", -- $0cd6d
          52590 => x"00", -- $0cd6e
          52591 => x"00", -- $0cd6f
          52592 => x"00", -- $0cd70
          52593 => x"00", -- $0cd71
          52594 => x"00", -- $0cd72
          52595 => x"00", -- $0cd73
          52596 => x"00", -- $0cd74
          52597 => x"00", -- $0cd75
          52598 => x"00", -- $0cd76
          52599 => x"00", -- $0cd77
          52600 => x"00", -- $0cd78
          52601 => x"00", -- $0cd79
          52602 => x"00", -- $0cd7a
          52603 => x"00", -- $0cd7b
          52604 => x"00", -- $0cd7c
          52605 => x"00", -- $0cd7d
          52606 => x"00", -- $0cd7e
          52607 => x"00", -- $0cd7f
          52608 => x"00", -- $0cd80
          52609 => x"00", -- $0cd81
          52610 => x"00", -- $0cd82
          52611 => x"00", -- $0cd83
          52612 => x"00", -- $0cd84
          52613 => x"00", -- $0cd85
          52614 => x"00", -- $0cd86
          52615 => x"00", -- $0cd87
          52616 => x"00", -- $0cd88
          52617 => x"00", -- $0cd89
          52618 => x"00", -- $0cd8a
          52619 => x"00", -- $0cd8b
          52620 => x"00", -- $0cd8c
          52621 => x"00", -- $0cd8d
          52622 => x"00", -- $0cd8e
          52623 => x"00", -- $0cd8f
          52624 => x"00", -- $0cd90
          52625 => x"00", -- $0cd91
          52626 => x"00", -- $0cd92
          52627 => x"00", -- $0cd93
          52628 => x"00", -- $0cd94
          52629 => x"00", -- $0cd95
          52630 => x"00", -- $0cd96
          52631 => x"00", -- $0cd97
          52632 => x"00", -- $0cd98
          52633 => x"00", -- $0cd99
          52634 => x"00", -- $0cd9a
          52635 => x"00", -- $0cd9b
          52636 => x"00", -- $0cd9c
          52637 => x"00", -- $0cd9d
          52638 => x"00", -- $0cd9e
          52639 => x"00", -- $0cd9f
          52640 => x"00", -- $0cda0
          52641 => x"00", -- $0cda1
          52642 => x"00", -- $0cda2
          52643 => x"00", -- $0cda3
          52644 => x"00", -- $0cda4
          52645 => x"00", -- $0cda5
          52646 => x"00", -- $0cda6
          52647 => x"00", -- $0cda7
          52648 => x"00", -- $0cda8
          52649 => x"00", -- $0cda9
          52650 => x"00", -- $0cdaa
          52651 => x"00", -- $0cdab
          52652 => x"00", -- $0cdac
          52653 => x"00", -- $0cdad
          52654 => x"00", -- $0cdae
          52655 => x"00", -- $0cdaf
          52656 => x"00", -- $0cdb0
          52657 => x"00", -- $0cdb1
          52658 => x"00", -- $0cdb2
          52659 => x"00", -- $0cdb3
          52660 => x"00", -- $0cdb4
          52661 => x"00", -- $0cdb5
          52662 => x"00", -- $0cdb6
          52663 => x"00", -- $0cdb7
          52664 => x"00", -- $0cdb8
          52665 => x"00", -- $0cdb9
          52666 => x"00", -- $0cdba
          52667 => x"00", -- $0cdbb
          52668 => x"00", -- $0cdbc
          52669 => x"00", -- $0cdbd
          52670 => x"00", -- $0cdbe
          52671 => x"00", -- $0cdbf
          52672 => x"00", -- $0cdc0
          52673 => x"00", -- $0cdc1
          52674 => x"00", -- $0cdc2
          52675 => x"00", -- $0cdc3
          52676 => x"00", -- $0cdc4
          52677 => x"00", -- $0cdc5
          52678 => x"00", -- $0cdc6
          52679 => x"00", -- $0cdc7
          52680 => x"00", -- $0cdc8
          52681 => x"00", -- $0cdc9
          52682 => x"00", -- $0cdca
          52683 => x"00", -- $0cdcb
          52684 => x"00", -- $0cdcc
          52685 => x"00", -- $0cdcd
          52686 => x"00", -- $0cdce
          52687 => x"00", -- $0cdcf
          52688 => x"00", -- $0cdd0
          52689 => x"00", -- $0cdd1
          52690 => x"00", -- $0cdd2
          52691 => x"00", -- $0cdd3
          52692 => x"00", -- $0cdd4
          52693 => x"00", -- $0cdd5
          52694 => x"00", -- $0cdd6
          52695 => x"00", -- $0cdd7
          52696 => x"00", -- $0cdd8
          52697 => x"00", -- $0cdd9
          52698 => x"00", -- $0cdda
          52699 => x"00", -- $0cddb
          52700 => x"00", -- $0cddc
          52701 => x"00", -- $0cddd
          52702 => x"00", -- $0cdde
          52703 => x"00", -- $0cddf
          52704 => x"00", -- $0cde0
          52705 => x"00", -- $0cde1
          52706 => x"00", -- $0cde2
          52707 => x"00", -- $0cde3
          52708 => x"00", -- $0cde4
          52709 => x"00", -- $0cde5
          52710 => x"00", -- $0cde6
          52711 => x"00", -- $0cde7
          52712 => x"00", -- $0cde8
          52713 => x"00", -- $0cde9
          52714 => x"00", -- $0cdea
          52715 => x"00", -- $0cdeb
          52716 => x"00", -- $0cdec
          52717 => x"00", -- $0cded
          52718 => x"00", -- $0cdee
          52719 => x"00", -- $0cdef
          52720 => x"00", -- $0cdf0
          52721 => x"00", -- $0cdf1
          52722 => x"00", -- $0cdf2
          52723 => x"00", -- $0cdf3
          52724 => x"00", -- $0cdf4
          52725 => x"00", -- $0cdf5
          52726 => x"00", -- $0cdf6
          52727 => x"00", -- $0cdf7
          52728 => x"00", -- $0cdf8
          52729 => x"00", -- $0cdf9
          52730 => x"00", -- $0cdfa
          52731 => x"00", -- $0cdfb
          52732 => x"00", -- $0cdfc
          52733 => x"00", -- $0cdfd
          52734 => x"00", -- $0cdfe
          52735 => x"00", -- $0cdff
          52736 => x"00", -- $0ce00
          52737 => x"00", -- $0ce01
          52738 => x"00", -- $0ce02
          52739 => x"00", -- $0ce03
          52740 => x"00", -- $0ce04
          52741 => x"00", -- $0ce05
          52742 => x"00", -- $0ce06
          52743 => x"00", -- $0ce07
          52744 => x"00", -- $0ce08
          52745 => x"00", -- $0ce09
          52746 => x"00", -- $0ce0a
          52747 => x"00", -- $0ce0b
          52748 => x"00", -- $0ce0c
          52749 => x"00", -- $0ce0d
          52750 => x"00", -- $0ce0e
          52751 => x"00", -- $0ce0f
          52752 => x"00", -- $0ce10
          52753 => x"00", -- $0ce11
          52754 => x"00", -- $0ce12
          52755 => x"00", -- $0ce13
          52756 => x"00", -- $0ce14
          52757 => x"00", -- $0ce15
          52758 => x"00", -- $0ce16
          52759 => x"00", -- $0ce17
          52760 => x"00", -- $0ce18
          52761 => x"00", -- $0ce19
          52762 => x"00", -- $0ce1a
          52763 => x"00", -- $0ce1b
          52764 => x"00", -- $0ce1c
          52765 => x"00", -- $0ce1d
          52766 => x"00", -- $0ce1e
          52767 => x"00", -- $0ce1f
          52768 => x"00", -- $0ce20
          52769 => x"00", -- $0ce21
          52770 => x"00", -- $0ce22
          52771 => x"00", -- $0ce23
          52772 => x"00", -- $0ce24
          52773 => x"00", -- $0ce25
          52774 => x"00", -- $0ce26
          52775 => x"00", -- $0ce27
          52776 => x"00", -- $0ce28
          52777 => x"00", -- $0ce29
          52778 => x"00", -- $0ce2a
          52779 => x"00", -- $0ce2b
          52780 => x"00", -- $0ce2c
          52781 => x"00", -- $0ce2d
          52782 => x"00", -- $0ce2e
          52783 => x"00", -- $0ce2f
          52784 => x"00", -- $0ce30
          52785 => x"00", -- $0ce31
          52786 => x"00", -- $0ce32
          52787 => x"00", -- $0ce33
          52788 => x"00", -- $0ce34
          52789 => x"00", -- $0ce35
          52790 => x"00", -- $0ce36
          52791 => x"00", -- $0ce37
          52792 => x"00", -- $0ce38
          52793 => x"00", -- $0ce39
          52794 => x"00", -- $0ce3a
          52795 => x"00", -- $0ce3b
          52796 => x"00", -- $0ce3c
          52797 => x"00", -- $0ce3d
          52798 => x"00", -- $0ce3e
          52799 => x"00", -- $0ce3f
          52800 => x"00", -- $0ce40
          52801 => x"00", -- $0ce41
          52802 => x"00", -- $0ce42
          52803 => x"00", -- $0ce43
          52804 => x"00", -- $0ce44
          52805 => x"00", -- $0ce45
          52806 => x"00", -- $0ce46
          52807 => x"00", -- $0ce47
          52808 => x"00", -- $0ce48
          52809 => x"00", -- $0ce49
          52810 => x"00", -- $0ce4a
          52811 => x"00", -- $0ce4b
          52812 => x"00", -- $0ce4c
          52813 => x"00", -- $0ce4d
          52814 => x"00", -- $0ce4e
          52815 => x"00", -- $0ce4f
          52816 => x"00", -- $0ce50
          52817 => x"00", -- $0ce51
          52818 => x"00", -- $0ce52
          52819 => x"00", -- $0ce53
          52820 => x"00", -- $0ce54
          52821 => x"00", -- $0ce55
          52822 => x"00", -- $0ce56
          52823 => x"00", -- $0ce57
          52824 => x"00", -- $0ce58
          52825 => x"00", -- $0ce59
          52826 => x"00", -- $0ce5a
          52827 => x"00", -- $0ce5b
          52828 => x"00", -- $0ce5c
          52829 => x"00", -- $0ce5d
          52830 => x"00", -- $0ce5e
          52831 => x"00", -- $0ce5f
          52832 => x"00", -- $0ce60
          52833 => x"00", -- $0ce61
          52834 => x"00", -- $0ce62
          52835 => x"00", -- $0ce63
          52836 => x"00", -- $0ce64
          52837 => x"00", -- $0ce65
          52838 => x"00", -- $0ce66
          52839 => x"00", -- $0ce67
          52840 => x"00", -- $0ce68
          52841 => x"00", -- $0ce69
          52842 => x"00", -- $0ce6a
          52843 => x"00", -- $0ce6b
          52844 => x"00", -- $0ce6c
          52845 => x"00", -- $0ce6d
          52846 => x"00", -- $0ce6e
          52847 => x"00", -- $0ce6f
          52848 => x"00", -- $0ce70
          52849 => x"00", -- $0ce71
          52850 => x"00", -- $0ce72
          52851 => x"00", -- $0ce73
          52852 => x"00", -- $0ce74
          52853 => x"00", -- $0ce75
          52854 => x"00", -- $0ce76
          52855 => x"00", -- $0ce77
          52856 => x"00", -- $0ce78
          52857 => x"00", -- $0ce79
          52858 => x"00", -- $0ce7a
          52859 => x"00", -- $0ce7b
          52860 => x"00", -- $0ce7c
          52861 => x"00", -- $0ce7d
          52862 => x"00", -- $0ce7e
          52863 => x"00", -- $0ce7f
          52864 => x"00", -- $0ce80
          52865 => x"00", -- $0ce81
          52866 => x"00", -- $0ce82
          52867 => x"00", -- $0ce83
          52868 => x"00", -- $0ce84
          52869 => x"00", -- $0ce85
          52870 => x"00", -- $0ce86
          52871 => x"00", -- $0ce87
          52872 => x"00", -- $0ce88
          52873 => x"00", -- $0ce89
          52874 => x"00", -- $0ce8a
          52875 => x"00", -- $0ce8b
          52876 => x"00", -- $0ce8c
          52877 => x"00", -- $0ce8d
          52878 => x"00", -- $0ce8e
          52879 => x"00", -- $0ce8f
          52880 => x"00", -- $0ce90
          52881 => x"00", -- $0ce91
          52882 => x"00", -- $0ce92
          52883 => x"00", -- $0ce93
          52884 => x"00", -- $0ce94
          52885 => x"00", -- $0ce95
          52886 => x"00", -- $0ce96
          52887 => x"00", -- $0ce97
          52888 => x"00", -- $0ce98
          52889 => x"00", -- $0ce99
          52890 => x"00", -- $0ce9a
          52891 => x"00", -- $0ce9b
          52892 => x"00", -- $0ce9c
          52893 => x"00", -- $0ce9d
          52894 => x"00", -- $0ce9e
          52895 => x"00", -- $0ce9f
          52896 => x"00", -- $0cea0
          52897 => x"00", -- $0cea1
          52898 => x"00", -- $0cea2
          52899 => x"00", -- $0cea3
          52900 => x"00", -- $0cea4
          52901 => x"00", -- $0cea5
          52902 => x"00", -- $0cea6
          52903 => x"00", -- $0cea7
          52904 => x"00", -- $0cea8
          52905 => x"00", -- $0cea9
          52906 => x"00", -- $0ceaa
          52907 => x"00", -- $0ceab
          52908 => x"00", -- $0ceac
          52909 => x"00", -- $0cead
          52910 => x"00", -- $0ceae
          52911 => x"00", -- $0ceaf
          52912 => x"00", -- $0ceb0
          52913 => x"00", -- $0ceb1
          52914 => x"00", -- $0ceb2
          52915 => x"00", -- $0ceb3
          52916 => x"00", -- $0ceb4
          52917 => x"00", -- $0ceb5
          52918 => x"00", -- $0ceb6
          52919 => x"00", -- $0ceb7
          52920 => x"00", -- $0ceb8
          52921 => x"00", -- $0ceb9
          52922 => x"00", -- $0ceba
          52923 => x"00", -- $0cebb
          52924 => x"00", -- $0cebc
          52925 => x"00", -- $0cebd
          52926 => x"00", -- $0cebe
          52927 => x"00", -- $0cebf
          52928 => x"00", -- $0cec0
          52929 => x"00", -- $0cec1
          52930 => x"00", -- $0cec2
          52931 => x"00", -- $0cec3
          52932 => x"00", -- $0cec4
          52933 => x"00", -- $0cec5
          52934 => x"00", -- $0cec6
          52935 => x"00", -- $0cec7
          52936 => x"00", -- $0cec8
          52937 => x"00", -- $0cec9
          52938 => x"00", -- $0ceca
          52939 => x"00", -- $0cecb
          52940 => x"00", -- $0cecc
          52941 => x"00", -- $0cecd
          52942 => x"00", -- $0cece
          52943 => x"00", -- $0cecf
          52944 => x"00", -- $0ced0
          52945 => x"00", -- $0ced1
          52946 => x"00", -- $0ced2
          52947 => x"00", -- $0ced3
          52948 => x"00", -- $0ced4
          52949 => x"00", -- $0ced5
          52950 => x"00", -- $0ced6
          52951 => x"00", -- $0ced7
          52952 => x"00", -- $0ced8
          52953 => x"00", -- $0ced9
          52954 => x"00", -- $0ceda
          52955 => x"00", -- $0cedb
          52956 => x"00", -- $0cedc
          52957 => x"00", -- $0cedd
          52958 => x"00", -- $0cede
          52959 => x"00", -- $0cedf
          52960 => x"00", -- $0cee0
          52961 => x"00", -- $0cee1
          52962 => x"00", -- $0cee2
          52963 => x"00", -- $0cee3
          52964 => x"00", -- $0cee4
          52965 => x"00", -- $0cee5
          52966 => x"00", -- $0cee6
          52967 => x"00", -- $0cee7
          52968 => x"00", -- $0cee8
          52969 => x"00", -- $0cee9
          52970 => x"00", -- $0ceea
          52971 => x"00", -- $0ceeb
          52972 => x"00", -- $0ceec
          52973 => x"00", -- $0ceed
          52974 => x"00", -- $0ceee
          52975 => x"00", -- $0ceef
          52976 => x"00", -- $0cef0
          52977 => x"00", -- $0cef1
          52978 => x"00", -- $0cef2
          52979 => x"00", -- $0cef3
          52980 => x"00", -- $0cef4
          52981 => x"00", -- $0cef5
          52982 => x"00", -- $0cef6
          52983 => x"00", -- $0cef7
          52984 => x"00", -- $0cef8
          52985 => x"00", -- $0cef9
          52986 => x"00", -- $0cefa
          52987 => x"00", -- $0cefb
          52988 => x"00", -- $0cefc
          52989 => x"00", -- $0cefd
          52990 => x"00", -- $0cefe
          52991 => x"00", -- $0ceff
          52992 => x"00", -- $0cf00
          52993 => x"00", -- $0cf01
          52994 => x"00", -- $0cf02
          52995 => x"00", -- $0cf03
          52996 => x"00", -- $0cf04
          52997 => x"00", -- $0cf05
          52998 => x"00", -- $0cf06
          52999 => x"00", -- $0cf07
          53000 => x"00", -- $0cf08
          53001 => x"00", -- $0cf09
          53002 => x"00", -- $0cf0a
          53003 => x"00", -- $0cf0b
          53004 => x"00", -- $0cf0c
          53005 => x"00", -- $0cf0d
          53006 => x"00", -- $0cf0e
          53007 => x"00", -- $0cf0f
          53008 => x"00", -- $0cf10
          53009 => x"00", -- $0cf11
          53010 => x"00", -- $0cf12
          53011 => x"00", -- $0cf13
          53012 => x"00", -- $0cf14
          53013 => x"00", -- $0cf15
          53014 => x"00", -- $0cf16
          53015 => x"00", -- $0cf17
          53016 => x"00", -- $0cf18
          53017 => x"00", -- $0cf19
          53018 => x"00", -- $0cf1a
          53019 => x"00", -- $0cf1b
          53020 => x"00", -- $0cf1c
          53021 => x"00", -- $0cf1d
          53022 => x"00", -- $0cf1e
          53023 => x"00", -- $0cf1f
          53024 => x"00", -- $0cf20
          53025 => x"00", -- $0cf21
          53026 => x"00", -- $0cf22
          53027 => x"00", -- $0cf23
          53028 => x"00", -- $0cf24
          53029 => x"00", -- $0cf25
          53030 => x"00", -- $0cf26
          53031 => x"00", -- $0cf27
          53032 => x"00", -- $0cf28
          53033 => x"00", -- $0cf29
          53034 => x"00", -- $0cf2a
          53035 => x"00", -- $0cf2b
          53036 => x"00", -- $0cf2c
          53037 => x"00", -- $0cf2d
          53038 => x"00", -- $0cf2e
          53039 => x"00", -- $0cf2f
          53040 => x"00", -- $0cf30
          53041 => x"00", -- $0cf31
          53042 => x"00", -- $0cf32
          53043 => x"00", -- $0cf33
          53044 => x"00", -- $0cf34
          53045 => x"00", -- $0cf35
          53046 => x"00", -- $0cf36
          53047 => x"00", -- $0cf37
          53048 => x"00", -- $0cf38
          53049 => x"00", -- $0cf39
          53050 => x"00", -- $0cf3a
          53051 => x"00", -- $0cf3b
          53052 => x"00", -- $0cf3c
          53053 => x"00", -- $0cf3d
          53054 => x"00", -- $0cf3e
          53055 => x"00", -- $0cf3f
          53056 => x"00", -- $0cf40
          53057 => x"00", -- $0cf41
          53058 => x"00", -- $0cf42
          53059 => x"00", -- $0cf43
          53060 => x"00", -- $0cf44
          53061 => x"00", -- $0cf45
          53062 => x"00", -- $0cf46
          53063 => x"00", -- $0cf47
          53064 => x"00", -- $0cf48
          53065 => x"00", -- $0cf49
          53066 => x"00", -- $0cf4a
          53067 => x"00", -- $0cf4b
          53068 => x"00", -- $0cf4c
          53069 => x"00", -- $0cf4d
          53070 => x"00", -- $0cf4e
          53071 => x"00", -- $0cf4f
          53072 => x"00", -- $0cf50
          53073 => x"00", -- $0cf51
          53074 => x"00", -- $0cf52
          53075 => x"00", -- $0cf53
          53076 => x"00", -- $0cf54
          53077 => x"00", -- $0cf55
          53078 => x"00", -- $0cf56
          53079 => x"00", -- $0cf57
          53080 => x"00", -- $0cf58
          53081 => x"00", -- $0cf59
          53082 => x"00", -- $0cf5a
          53083 => x"00", -- $0cf5b
          53084 => x"00", -- $0cf5c
          53085 => x"00", -- $0cf5d
          53086 => x"00", -- $0cf5e
          53087 => x"00", -- $0cf5f
          53088 => x"00", -- $0cf60
          53089 => x"00", -- $0cf61
          53090 => x"00", -- $0cf62
          53091 => x"00", -- $0cf63
          53092 => x"00", -- $0cf64
          53093 => x"00", -- $0cf65
          53094 => x"00", -- $0cf66
          53095 => x"00", -- $0cf67
          53096 => x"00", -- $0cf68
          53097 => x"00", -- $0cf69
          53098 => x"00", -- $0cf6a
          53099 => x"00", -- $0cf6b
          53100 => x"00", -- $0cf6c
          53101 => x"00", -- $0cf6d
          53102 => x"00", -- $0cf6e
          53103 => x"00", -- $0cf6f
          53104 => x"00", -- $0cf70
          53105 => x"00", -- $0cf71
          53106 => x"00", -- $0cf72
          53107 => x"00", -- $0cf73
          53108 => x"00", -- $0cf74
          53109 => x"00", -- $0cf75
          53110 => x"00", -- $0cf76
          53111 => x"00", -- $0cf77
          53112 => x"00", -- $0cf78
          53113 => x"00", -- $0cf79
          53114 => x"00", -- $0cf7a
          53115 => x"00", -- $0cf7b
          53116 => x"00", -- $0cf7c
          53117 => x"00", -- $0cf7d
          53118 => x"00", -- $0cf7e
          53119 => x"00", -- $0cf7f
          53120 => x"00", -- $0cf80
          53121 => x"00", -- $0cf81
          53122 => x"00", -- $0cf82
          53123 => x"00", -- $0cf83
          53124 => x"00", -- $0cf84
          53125 => x"00", -- $0cf85
          53126 => x"00", -- $0cf86
          53127 => x"00", -- $0cf87
          53128 => x"00", -- $0cf88
          53129 => x"00", -- $0cf89
          53130 => x"00", -- $0cf8a
          53131 => x"00", -- $0cf8b
          53132 => x"00", -- $0cf8c
          53133 => x"00", -- $0cf8d
          53134 => x"00", -- $0cf8e
          53135 => x"00", -- $0cf8f
          53136 => x"00", -- $0cf90
          53137 => x"00", -- $0cf91
          53138 => x"00", -- $0cf92
          53139 => x"00", -- $0cf93
          53140 => x"00", -- $0cf94
          53141 => x"00", -- $0cf95
          53142 => x"00", -- $0cf96
          53143 => x"00", -- $0cf97
          53144 => x"00", -- $0cf98
          53145 => x"00", -- $0cf99
          53146 => x"00", -- $0cf9a
          53147 => x"00", -- $0cf9b
          53148 => x"00", -- $0cf9c
          53149 => x"00", -- $0cf9d
          53150 => x"00", -- $0cf9e
          53151 => x"00", -- $0cf9f
          53152 => x"00", -- $0cfa0
          53153 => x"00", -- $0cfa1
          53154 => x"00", -- $0cfa2
          53155 => x"00", -- $0cfa3
          53156 => x"00", -- $0cfa4
          53157 => x"00", -- $0cfa5
          53158 => x"00", -- $0cfa6
          53159 => x"00", -- $0cfa7
          53160 => x"00", -- $0cfa8
          53161 => x"00", -- $0cfa9
          53162 => x"00", -- $0cfaa
          53163 => x"00", -- $0cfab
          53164 => x"00", -- $0cfac
          53165 => x"00", -- $0cfad
          53166 => x"00", -- $0cfae
          53167 => x"00", -- $0cfaf
          53168 => x"00", -- $0cfb0
          53169 => x"00", -- $0cfb1
          53170 => x"00", -- $0cfb2
          53171 => x"00", -- $0cfb3
          53172 => x"00", -- $0cfb4
          53173 => x"00", -- $0cfb5
          53174 => x"00", -- $0cfb6
          53175 => x"00", -- $0cfb7
          53176 => x"00", -- $0cfb8
          53177 => x"00", -- $0cfb9
          53178 => x"00", -- $0cfba
          53179 => x"00", -- $0cfbb
          53180 => x"00", -- $0cfbc
          53181 => x"00", -- $0cfbd
          53182 => x"00", -- $0cfbe
          53183 => x"00", -- $0cfbf
          53184 => x"00", -- $0cfc0
          53185 => x"00", -- $0cfc1
          53186 => x"00", -- $0cfc2
          53187 => x"00", -- $0cfc3
          53188 => x"00", -- $0cfc4
          53189 => x"00", -- $0cfc5
          53190 => x"00", -- $0cfc6
          53191 => x"00", -- $0cfc7
          53192 => x"00", -- $0cfc8
          53193 => x"00", -- $0cfc9
          53194 => x"00", -- $0cfca
          53195 => x"00", -- $0cfcb
          53196 => x"00", -- $0cfcc
          53197 => x"00", -- $0cfcd
          53198 => x"00", -- $0cfce
          53199 => x"00", -- $0cfcf
          53200 => x"00", -- $0cfd0
          53201 => x"00", -- $0cfd1
          53202 => x"00", -- $0cfd2
          53203 => x"00", -- $0cfd3
          53204 => x"00", -- $0cfd4
          53205 => x"00", -- $0cfd5
          53206 => x"00", -- $0cfd6
          53207 => x"00", -- $0cfd7
          53208 => x"00", -- $0cfd8
          53209 => x"00", -- $0cfd9
          53210 => x"00", -- $0cfda
          53211 => x"00", -- $0cfdb
          53212 => x"00", -- $0cfdc
          53213 => x"00", -- $0cfdd
          53214 => x"00", -- $0cfde
          53215 => x"00", -- $0cfdf
          53216 => x"00", -- $0cfe0
          53217 => x"00", -- $0cfe1
          53218 => x"00", -- $0cfe2
          53219 => x"00", -- $0cfe3
          53220 => x"00", -- $0cfe4
          53221 => x"00", -- $0cfe5
          53222 => x"00", -- $0cfe6
          53223 => x"00", -- $0cfe7
          53224 => x"00", -- $0cfe8
          53225 => x"00", -- $0cfe9
          53226 => x"00", -- $0cfea
          53227 => x"00", -- $0cfeb
          53228 => x"00", -- $0cfec
          53229 => x"00", -- $0cfed
          53230 => x"00", -- $0cfee
          53231 => x"00", -- $0cfef
          53232 => x"00", -- $0cff0
          53233 => x"00", -- $0cff1
          53234 => x"00", -- $0cff2
          53235 => x"00", -- $0cff3
          53236 => x"00", -- $0cff4
          53237 => x"00", -- $0cff5
          53238 => x"00", -- $0cff6
          53239 => x"00", -- $0cff7
          53240 => x"00", -- $0cff8
          53241 => x"00", -- $0cff9
          53242 => x"00", -- $0cffa
          53243 => x"00", -- $0cffb
          53244 => x"00", -- $0cffc
          53245 => x"00", -- $0cffd
          53246 => x"00", -- $0cffe
          53247 => x"00", -- $0cfff
          53248 => x"00", -- $0d000
          53249 => x"00", -- $0d001
          53250 => x"00", -- $0d002
          53251 => x"00", -- $0d003
          53252 => x"00", -- $0d004
          53253 => x"00", -- $0d005
          53254 => x"00", -- $0d006
          53255 => x"00", -- $0d007
          53256 => x"00", -- $0d008
          53257 => x"00", -- $0d009
          53258 => x"00", -- $0d00a
          53259 => x"00", -- $0d00b
          53260 => x"00", -- $0d00c
          53261 => x"00", -- $0d00d
          53262 => x"00", -- $0d00e
          53263 => x"00", -- $0d00f
          53264 => x"00", -- $0d010
          53265 => x"00", -- $0d011
          53266 => x"00", -- $0d012
          53267 => x"00", -- $0d013
          53268 => x"00", -- $0d014
          53269 => x"00", -- $0d015
          53270 => x"00", -- $0d016
          53271 => x"00", -- $0d017
          53272 => x"00", -- $0d018
          53273 => x"00", -- $0d019
          53274 => x"00", -- $0d01a
          53275 => x"00", -- $0d01b
          53276 => x"00", -- $0d01c
          53277 => x"00", -- $0d01d
          53278 => x"00", -- $0d01e
          53279 => x"00", -- $0d01f
          53280 => x"00", -- $0d020
          53281 => x"00", -- $0d021
          53282 => x"00", -- $0d022
          53283 => x"00", -- $0d023
          53284 => x"00", -- $0d024
          53285 => x"00", -- $0d025
          53286 => x"00", -- $0d026
          53287 => x"00", -- $0d027
          53288 => x"00", -- $0d028
          53289 => x"00", -- $0d029
          53290 => x"00", -- $0d02a
          53291 => x"00", -- $0d02b
          53292 => x"00", -- $0d02c
          53293 => x"00", -- $0d02d
          53294 => x"00", -- $0d02e
          53295 => x"00", -- $0d02f
          53296 => x"00", -- $0d030
          53297 => x"00", -- $0d031
          53298 => x"00", -- $0d032
          53299 => x"00", -- $0d033
          53300 => x"00", -- $0d034
          53301 => x"00", -- $0d035
          53302 => x"00", -- $0d036
          53303 => x"00", -- $0d037
          53304 => x"00", -- $0d038
          53305 => x"00", -- $0d039
          53306 => x"00", -- $0d03a
          53307 => x"00", -- $0d03b
          53308 => x"00", -- $0d03c
          53309 => x"00", -- $0d03d
          53310 => x"00", -- $0d03e
          53311 => x"00", -- $0d03f
          53312 => x"00", -- $0d040
          53313 => x"00", -- $0d041
          53314 => x"00", -- $0d042
          53315 => x"00", -- $0d043
          53316 => x"00", -- $0d044
          53317 => x"00", -- $0d045
          53318 => x"00", -- $0d046
          53319 => x"00", -- $0d047
          53320 => x"00", -- $0d048
          53321 => x"00", -- $0d049
          53322 => x"00", -- $0d04a
          53323 => x"00", -- $0d04b
          53324 => x"00", -- $0d04c
          53325 => x"00", -- $0d04d
          53326 => x"00", -- $0d04e
          53327 => x"00", -- $0d04f
          53328 => x"00", -- $0d050
          53329 => x"00", -- $0d051
          53330 => x"00", -- $0d052
          53331 => x"00", -- $0d053
          53332 => x"00", -- $0d054
          53333 => x"00", -- $0d055
          53334 => x"00", -- $0d056
          53335 => x"00", -- $0d057
          53336 => x"00", -- $0d058
          53337 => x"00", -- $0d059
          53338 => x"00", -- $0d05a
          53339 => x"00", -- $0d05b
          53340 => x"00", -- $0d05c
          53341 => x"00", -- $0d05d
          53342 => x"00", -- $0d05e
          53343 => x"00", -- $0d05f
          53344 => x"00", -- $0d060
          53345 => x"00", -- $0d061
          53346 => x"00", -- $0d062
          53347 => x"00", -- $0d063
          53348 => x"00", -- $0d064
          53349 => x"00", -- $0d065
          53350 => x"00", -- $0d066
          53351 => x"00", -- $0d067
          53352 => x"00", -- $0d068
          53353 => x"00", -- $0d069
          53354 => x"00", -- $0d06a
          53355 => x"00", -- $0d06b
          53356 => x"00", -- $0d06c
          53357 => x"00", -- $0d06d
          53358 => x"00", -- $0d06e
          53359 => x"00", -- $0d06f
          53360 => x"00", -- $0d070
          53361 => x"00", -- $0d071
          53362 => x"00", -- $0d072
          53363 => x"00", -- $0d073
          53364 => x"00", -- $0d074
          53365 => x"00", -- $0d075
          53366 => x"00", -- $0d076
          53367 => x"00", -- $0d077
          53368 => x"00", -- $0d078
          53369 => x"00", -- $0d079
          53370 => x"00", -- $0d07a
          53371 => x"00", -- $0d07b
          53372 => x"00", -- $0d07c
          53373 => x"00", -- $0d07d
          53374 => x"00", -- $0d07e
          53375 => x"00", -- $0d07f
          53376 => x"00", -- $0d080
          53377 => x"00", -- $0d081
          53378 => x"00", -- $0d082
          53379 => x"00", -- $0d083
          53380 => x"00", -- $0d084
          53381 => x"00", -- $0d085
          53382 => x"00", -- $0d086
          53383 => x"00", -- $0d087
          53384 => x"00", -- $0d088
          53385 => x"00", -- $0d089
          53386 => x"00", -- $0d08a
          53387 => x"00", -- $0d08b
          53388 => x"00", -- $0d08c
          53389 => x"00", -- $0d08d
          53390 => x"00", -- $0d08e
          53391 => x"00", -- $0d08f
          53392 => x"00", -- $0d090
          53393 => x"00", -- $0d091
          53394 => x"00", -- $0d092
          53395 => x"00", -- $0d093
          53396 => x"00", -- $0d094
          53397 => x"00", -- $0d095
          53398 => x"00", -- $0d096
          53399 => x"00", -- $0d097
          53400 => x"00", -- $0d098
          53401 => x"00", -- $0d099
          53402 => x"00", -- $0d09a
          53403 => x"00", -- $0d09b
          53404 => x"00", -- $0d09c
          53405 => x"00", -- $0d09d
          53406 => x"00", -- $0d09e
          53407 => x"00", -- $0d09f
          53408 => x"00", -- $0d0a0
          53409 => x"00", -- $0d0a1
          53410 => x"00", -- $0d0a2
          53411 => x"00", -- $0d0a3
          53412 => x"00", -- $0d0a4
          53413 => x"00", -- $0d0a5
          53414 => x"00", -- $0d0a6
          53415 => x"00", -- $0d0a7
          53416 => x"00", -- $0d0a8
          53417 => x"00", -- $0d0a9
          53418 => x"00", -- $0d0aa
          53419 => x"00", -- $0d0ab
          53420 => x"00", -- $0d0ac
          53421 => x"00", -- $0d0ad
          53422 => x"00", -- $0d0ae
          53423 => x"00", -- $0d0af
          53424 => x"00", -- $0d0b0
          53425 => x"00", -- $0d0b1
          53426 => x"00", -- $0d0b2
          53427 => x"00", -- $0d0b3
          53428 => x"00", -- $0d0b4
          53429 => x"00", -- $0d0b5
          53430 => x"00", -- $0d0b6
          53431 => x"00", -- $0d0b7
          53432 => x"00", -- $0d0b8
          53433 => x"00", -- $0d0b9
          53434 => x"00", -- $0d0ba
          53435 => x"00", -- $0d0bb
          53436 => x"00", -- $0d0bc
          53437 => x"00", -- $0d0bd
          53438 => x"00", -- $0d0be
          53439 => x"00", -- $0d0bf
          53440 => x"00", -- $0d0c0
          53441 => x"00", -- $0d0c1
          53442 => x"00", -- $0d0c2
          53443 => x"00", -- $0d0c3
          53444 => x"00", -- $0d0c4
          53445 => x"00", -- $0d0c5
          53446 => x"00", -- $0d0c6
          53447 => x"00", -- $0d0c7
          53448 => x"00", -- $0d0c8
          53449 => x"00", -- $0d0c9
          53450 => x"00", -- $0d0ca
          53451 => x"00", -- $0d0cb
          53452 => x"00", -- $0d0cc
          53453 => x"00", -- $0d0cd
          53454 => x"00", -- $0d0ce
          53455 => x"00", -- $0d0cf
          53456 => x"00", -- $0d0d0
          53457 => x"00", -- $0d0d1
          53458 => x"00", -- $0d0d2
          53459 => x"00", -- $0d0d3
          53460 => x"00", -- $0d0d4
          53461 => x"00", -- $0d0d5
          53462 => x"00", -- $0d0d6
          53463 => x"00", -- $0d0d7
          53464 => x"00", -- $0d0d8
          53465 => x"00", -- $0d0d9
          53466 => x"00", -- $0d0da
          53467 => x"00", -- $0d0db
          53468 => x"00", -- $0d0dc
          53469 => x"00", -- $0d0dd
          53470 => x"00", -- $0d0de
          53471 => x"00", -- $0d0df
          53472 => x"00", -- $0d0e0
          53473 => x"00", -- $0d0e1
          53474 => x"00", -- $0d0e2
          53475 => x"00", -- $0d0e3
          53476 => x"00", -- $0d0e4
          53477 => x"00", -- $0d0e5
          53478 => x"00", -- $0d0e6
          53479 => x"00", -- $0d0e7
          53480 => x"00", -- $0d0e8
          53481 => x"00", -- $0d0e9
          53482 => x"00", -- $0d0ea
          53483 => x"00", -- $0d0eb
          53484 => x"00", -- $0d0ec
          53485 => x"00", -- $0d0ed
          53486 => x"00", -- $0d0ee
          53487 => x"00", -- $0d0ef
          53488 => x"00", -- $0d0f0
          53489 => x"00", -- $0d0f1
          53490 => x"00", -- $0d0f2
          53491 => x"00", -- $0d0f3
          53492 => x"00", -- $0d0f4
          53493 => x"00", -- $0d0f5
          53494 => x"00", -- $0d0f6
          53495 => x"00", -- $0d0f7
          53496 => x"00", -- $0d0f8
          53497 => x"00", -- $0d0f9
          53498 => x"00", -- $0d0fa
          53499 => x"00", -- $0d0fb
          53500 => x"00", -- $0d0fc
          53501 => x"00", -- $0d0fd
          53502 => x"00", -- $0d0fe
          53503 => x"00", -- $0d0ff
          53504 => x"00", -- $0d100
          53505 => x"00", -- $0d101
          53506 => x"00", -- $0d102
          53507 => x"00", -- $0d103
          53508 => x"00", -- $0d104
          53509 => x"00", -- $0d105
          53510 => x"00", -- $0d106
          53511 => x"00", -- $0d107
          53512 => x"00", -- $0d108
          53513 => x"00", -- $0d109
          53514 => x"00", -- $0d10a
          53515 => x"00", -- $0d10b
          53516 => x"00", -- $0d10c
          53517 => x"00", -- $0d10d
          53518 => x"00", -- $0d10e
          53519 => x"00", -- $0d10f
          53520 => x"00", -- $0d110
          53521 => x"00", -- $0d111
          53522 => x"00", -- $0d112
          53523 => x"00", -- $0d113
          53524 => x"00", -- $0d114
          53525 => x"00", -- $0d115
          53526 => x"00", -- $0d116
          53527 => x"00", -- $0d117
          53528 => x"00", -- $0d118
          53529 => x"00", -- $0d119
          53530 => x"00", -- $0d11a
          53531 => x"00", -- $0d11b
          53532 => x"00", -- $0d11c
          53533 => x"00", -- $0d11d
          53534 => x"00", -- $0d11e
          53535 => x"00", -- $0d11f
          53536 => x"00", -- $0d120
          53537 => x"00", -- $0d121
          53538 => x"00", -- $0d122
          53539 => x"00", -- $0d123
          53540 => x"00", -- $0d124
          53541 => x"00", -- $0d125
          53542 => x"00", -- $0d126
          53543 => x"00", -- $0d127
          53544 => x"00", -- $0d128
          53545 => x"00", -- $0d129
          53546 => x"00", -- $0d12a
          53547 => x"00", -- $0d12b
          53548 => x"00", -- $0d12c
          53549 => x"00", -- $0d12d
          53550 => x"00", -- $0d12e
          53551 => x"00", -- $0d12f
          53552 => x"00", -- $0d130
          53553 => x"00", -- $0d131
          53554 => x"00", -- $0d132
          53555 => x"00", -- $0d133
          53556 => x"00", -- $0d134
          53557 => x"00", -- $0d135
          53558 => x"00", -- $0d136
          53559 => x"00", -- $0d137
          53560 => x"00", -- $0d138
          53561 => x"00", -- $0d139
          53562 => x"00", -- $0d13a
          53563 => x"00", -- $0d13b
          53564 => x"00", -- $0d13c
          53565 => x"00", -- $0d13d
          53566 => x"00", -- $0d13e
          53567 => x"00", -- $0d13f
          53568 => x"00", -- $0d140
          53569 => x"00", -- $0d141
          53570 => x"00", -- $0d142
          53571 => x"00", -- $0d143
          53572 => x"00", -- $0d144
          53573 => x"00", -- $0d145
          53574 => x"00", -- $0d146
          53575 => x"00", -- $0d147
          53576 => x"00", -- $0d148
          53577 => x"00", -- $0d149
          53578 => x"00", -- $0d14a
          53579 => x"00", -- $0d14b
          53580 => x"00", -- $0d14c
          53581 => x"00", -- $0d14d
          53582 => x"00", -- $0d14e
          53583 => x"00", -- $0d14f
          53584 => x"00", -- $0d150
          53585 => x"00", -- $0d151
          53586 => x"00", -- $0d152
          53587 => x"00", -- $0d153
          53588 => x"00", -- $0d154
          53589 => x"00", -- $0d155
          53590 => x"00", -- $0d156
          53591 => x"00", -- $0d157
          53592 => x"00", -- $0d158
          53593 => x"00", -- $0d159
          53594 => x"00", -- $0d15a
          53595 => x"00", -- $0d15b
          53596 => x"00", -- $0d15c
          53597 => x"00", -- $0d15d
          53598 => x"00", -- $0d15e
          53599 => x"00", -- $0d15f
          53600 => x"00", -- $0d160
          53601 => x"00", -- $0d161
          53602 => x"00", -- $0d162
          53603 => x"00", -- $0d163
          53604 => x"00", -- $0d164
          53605 => x"00", -- $0d165
          53606 => x"00", -- $0d166
          53607 => x"00", -- $0d167
          53608 => x"00", -- $0d168
          53609 => x"00", -- $0d169
          53610 => x"00", -- $0d16a
          53611 => x"00", -- $0d16b
          53612 => x"00", -- $0d16c
          53613 => x"00", -- $0d16d
          53614 => x"00", -- $0d16e
          53615 => x"00", -- $0d16f
          53616 => x"00", -- $0d170
          53617 => x"00", -- $0d171
          53618 => x"00", -- $0d172
          53619 => x"00", -- $0d173
          53620 => x"00", -- $0d174
          53621 => x"00", -- $0d175
          53622 => x"00", -- $0d176
          53623 => x"00", -- $0d177
          53624 => x"00", -- $0d178
          53625 => x"00", -- $0d179
          53626 => x"00", -- $0d17a
          53627 => x"00", -- $0d17b
          53628 => x"00", -- $0d17c
          53629 => x"00", -- $0d17d
          53630 => x"00", -- $0d17e
          53631 => x"00", -- $0d17f
          53632 => x"00", -- $0d180
          53633 => x"00", -- $0d181
          53634 => x"00", -- $0d182
          53635 => x"00", -- $0d183
          53636 => x"00", -- $0d184
          53637 => x"00", -- $0d185
          53638 => x"00", -- $0d186
          53639 => x"00", -- $0d187
          53640 => x"00", -- $0d188
          53641 => x"00", -- $0d189
          53642 => x"00", -- $0d18a
          53643 => x"00", -- $0d18b
          53644 => x"00", -- $0d18c
          53645 => x"00", -- $0d18d
          53646 => x"00", -- $0d18e
          53647 => x"00", -- $0d18f
          53648 => x"00", -- $0d190
          53649 => x"00", -- $0d191
          53650 => x"00", -- $0d192
          53651 => x"00", -- $0d193
          53652 => x"00", -- $0d194
          53653 => x"00", -- $0d195
          53654 => x"00", -- $0d196
          53655 => x"00", -- $0d197
          53656 => x"00", -- $0d198
          53657 => x"00", -- $0d199
          53658 => x"00", -- $0d19a
          53659 => x"00", -- $0d19b
          53660 => x"00", -- $0d19c
          53661 => x"00", -- $0d19d
          53662 => x"00", -- $0d19e
          53663 => x"00", -- $0d19f
          53664 => x"00", -- $0d1a0
          53665 => x"00", -- $0d1a1
          53666 => x"00", -- $0d1a2
          53667 => x"00", -- $0d1a3
          53668 => x"00", -- $0d1a4
          53669 => x"00", -- $0d1a5
          53670 => x"00", -- $0d1a6
          53671 => x"00", -- $0d1a7
          53672 => x"00", -- $0d1a8
          53673 => x"00", -- $0d1a9
          53674 => x"00", -- $0d1aa
          53675 => x"00", -- $0d1ab
          53676 => x"00", -- $0d1ac
          53677 => x"00", -- $0d1ad
          53678 => x"00", -- $0d1ae
          53679 => x"00", -- $0d1af
          53680 => x"00", -- $0d1b0
          53681 => x"00", -- $0d1b1
          53682 => x"00", -- $0d1b2
          53683 => x"00", -- $0d1b3
          53684 => x"00", -- $0d1b4
          53685 => x"00", -- $0d1b5
          53686 => x"00", -- $0d1b6
          53687 => x"00", -- $0d1b7
          53688 => x"00", -- $0d1b8
          53689 => x"00", -- $0d1b9
          53690 => x"00", -- $0d1ba
          53691 => x"00", -- $0d1bb
          53692 => x"00", -- $0d1bc
          53693 => x"00", -- $0d1bd
          53694 => x"00", -- $0d1be
          53695 => x"00", -- $0d1bf
          53696 => x"00", -- $0d1c0
          53697 => x"00", -- $0d1c1
          53698 => x"00", -- $0d1c2
          53699 => x"00", -- $0d1c3
          53700 => x"00", -- $0d1c4
          53701 => x"00", -- $0d1c5
          53702 => x"00", -- $0d1c6
          53703 => x"00", -- $0d1c7
          53704 => x"00", -- $0d1c8
          53705 => x"00", -- $0d1c9
          53706 => x"00", -- $0d1ca
          53707 => x"00", -- $0d1cb
          53708 => x"00", -- $0d1cc
          53709 => x"00", -- $0d1cd
          53710 => x"00", -- $0d1ce
          53711 => x"00", -- $0d1cf
          53712 => x"00", -- $0d1d0
          53713 => x"00", -- $0d1d1
          53714 => x"00", -- $0d1d2
          53715 => x"00", -- $0d1d3
          53716 => x"00", -- $0d1d4
          53717 => x"00", -- $0d1d5
          53718 => x"00", -- $0d1d6
          53719 => x"00", -- $0d1d7
          53720 => x"00", -- $0d1d8
          53721 => x"00", -- $0d1d9
          53722 => x"00", -- $0d1da
          53723 => x"00", -- $0d1db
          53724 => x"00", -- $0d1dc
          53725 => x"00", -- $0d1dd
          53726 => x"00", -- $0d1de
          53727 => x"00", -- $0d1df
          53728 => x"00", -- $0d1e0
          53729 => x"00", -- $0d1e1
          53730 => x"00", -- $0d1e2
          53731 => x"00", -- $0d1e3
          53732 => x"00", -- $0d1e4
          53733 => x"00", -- $0d1e5
          53734 => x"00", -- $0d1e6
          53735 => x"00", -- $0d1e7
          53736 => x"00", -- $0d1e8
          53737 => x"00", -- $0d1e9
          53738 => x"00", -- $0d1ea
          53739 => x"00", -- $0d1eb
          53740 => x"00", -- $0d1ec
          53741 => x"00", -- $0d1ed
          53742 => x"00", -- $0d1ee
          53743 => x"00", -- $0d1ef
          53744 => x"00", -- $0d1f0
          53745 => x"00", -- $0d1f1
          53746 => x"00", -- $0d1f2
          53747 => x"00", -- $0d1f3
          53748 => x"00", -- $0d1f4
          53749 => x"00", -- $0d1f5
          53750 => x"00", -- $0d1f6
          53751 => x"00", -- $0d1f7
          53752 => x"00", -- $0d1f8
          53753 => x"00", -- $0d1f9
          53754 => x"00", -- $0d1fa
          53755 => x"00", -- $0d1fb
          53756 => x"00", -- $0d1fc
          53757 => x"00", -- $0d1fd
          53758 => x"00", -- $0d1fe
          53759 => x"00", -- $0d1ff
          53760 => x"00", -- $0d200
          53761 => x"00", -- $0d201
          53762 => x"00", -- $0d202
          53763 => x"00", -- $0d203
          53764 => x"00", -- $0d204
          53765 => x"00", -- $0d205
          53766 => x"00", -- $0d206
          53767 => x"00", -- $0d207
          53768 => x"00", -- $0d208
          53769 => x"00", -- $0d209
          53770 => x"00", -- $0d20a
          53771 => x"00", -- $0d20b
          53772 => x"00", -- $0d20c
          53773 => x"00", -- $0d20d
          53774 => x"00", -- $0d20e
          53775 => x"00", -- $0d20f
          53776 => x"00", -- $0d210
          53777 => x"00", -- $0d211
          53778 => x"00", -- $0d212
          53779 => x"00", -- $0d213
          53780 => x"00", -- $0d214
          53781 => x"00", -- $0d215
          53782 => x"00", -- $0d216
          53783 => x"00", -- $0d217
          53784 => x"00", -- $0d218
          53785 => x"00", -- $0d219
          53786 => x"00", -- $0d21a
          53787 => x"00", -- $0d21b
          53788 => x"00", -- $0d21c
          53789 => x"00", -- $0d21d
          53790 => x"00", -- $0d21e
          53791 => x"00", -- $0d21f
          53792 => x"00", -- $0d220
          53793 => x"00", -- $0d221
          53794 => x"00", -- $0d222
          53795 => x"00", -- $0d223
          53796 => x"00", -- $0d224
          53797 => x"00", -- $0d225
          53798 => x"00", -- $0d226
          53799 => x"00", -- $0d227
          53800 => x"00", -- $0d228
          53801 => x"00", -- $0d229
          53802 => x"00", -- $0d22a
          53803 => x"00", -- $0d22b
          53804 => x"00", -- $0d22c
          53805 => x"00", -- $0d22d
          53806 => x"00", -- $0d22e
          53807 => x"00", -- $0d22f
          53808 => x"00", -- $0d230
          53809 => x"00", -- $0d231
          53810 => x"00", -- $0d232
          53811 => x"00", -- $0d233
          53812 => x"00", -- $0d234
          53813 => x"00", -- $0d235
          53814 => x"00", -- $0d236
          53815 => x"00", -- $0d237
          53816 => x"00", -- $0d238
          53817 => x"00", -- $0d239
          53818 => x"00", -- $0d23a
          53819 => x"00", -- $0d23b
          53820 => x"00", -- $0d23c
          53821 => x"00", -- $0d23d
          53822 => x"00", -- $0d23e
          53823 => x"00", -- $0d23f
          53824 => x"00", -- $0d240
          53825 => x"00", -- $0d241
          53826 => x"00", -- $0d242
          53827 => x"00", -- $0d243
          53828 => x"00", -- $0d244
          53829 => x"00", -- $0d245
          53830 => x"00", -- $0d246
          53831 => x"00", -- $0d247
          53832 => x"00", -- $0d248
          53833 => x"00", -- $0d249
          53834 => x"00", -- $0d24a
          53835 => x"00", -- $0d24b
          53836 => x"00", -- $0d24c
          53837 => x"00", -- $0d24d
          53838 => x"00", -- $0d24e
          53839 => x"00", -- $0d24f
          53840 => x"00", -- $0d250
          53841 => x"00", -- $0d251
          53842 => x"00", -- $0d252
          53843 => x"00", -- $0d253
          53844 => x"00", -- $0d254
          53845 => x"00", -- $0d255
          53846 => x"00", -- $0d256
          53847 => x"00", -- $0d257
          53848 => x"00", -- $0d258
          53849 => x"00", -- $0d259
          53850 => x"00", -- $0d25a
          53851 => x"00", -- $0d25b
          53852 => x"00", -- $0d25c
          53853 => x"00", -- $0d25d
          53854 => x"00", -- $0d25e
          53855 => x"00", -- $0d25f
          53856 => x"00", -- $0d260
          53857 => x"00", -- $0d261
          53858 => x"00", -- $0d262
          53859 => x"00", -- $0d263
          53860 => x"00", -- $0d264
          53861 => x"00", -- $0d265
          53862 => x"00", -- $0d266
          53863 => x"00", -- $0d267
          53864 => x"00", -- $0d268
          53865 => x"00", -- $0d269
          53866 => x"00", -- $0d26a
          53867 => x"00", -- $0d26b
          53868 => x"00", -- $0d26c
          53869 => x"00", -- $0d26d
          53870 => x"00", -- $0d26e
          53871 => x"00", -- $0d26f
          53872 => x"00", -- $0d270
          53873 => x"00", -- $0d271
          53874 => x"00", -- $0d272
          53875 => x"00", -- $0d273
          53876 => x"00", -- $0d274
          53877 => x"00", -- $0d275
          53878 => x"00", -- $0d276
          53879 => x"00", -- $0d277
          53880 => x"00", -- $0d278
          53881 => x"00", -- $0d279
          53882 => x"00", -- $0d27a
          53883 => x"00", -- $0d27b
          53884 => x"00", -- $0d27c
          53885 => x"00", -- $0d27d
          53886 => x"00", -- $0d27e
          53887 => x"00", -- $0d27f
          53888 => x"00", -- $0d280
          53889 => x"00", -- $0d281
          53890 => x"00", -- $0d282
          53891 => x"00", -- $0d283
          53892 => x"00", -- $0d284
          53893 => x"00", -- $0d285
          53894 => x"00", -- $0d286
          53895 => x"00", -- $0d287
          53896 => x"00", -- $0d288
          53897 => x"00", -- $0d289
          53898 => x"00", -- $0d28a
          53899 => x"00", -- $0d28b
          53900 => x"00", -- $0d28c
          53901 => x"00", -- $0d28d
          53902 => x"00", -- $0d28e
          53903 => x"00", -- $0d28f
          53904 => x"00", -- $0d290
          53905 => x"00", -- $0d291
          53906 => x"00", -- $0d292
          53907 => x"00", -- $0d293
          53908 => x"00", -- $0d294
          53909 => x"00", -- $0d295
          53910 => x"00", -- $0d296
          53911 => x"00", -- $0d297
          53912 => x"00", -- $0d298
          53913 => x"00", -- $0d299
          53914 => x"00", -- $0d29a
          53915 => x"00", -- $0d29b
          53916 => x"00", -- $0d29c
          53917 => x"00", -- $0d29d
          53918 => x"00", -- $0d29e
          53919 => x"00", -- $0d29f
          53920 => x"00", -- $0d2a0
          53921 => x"00", -- $0d2a1
          53922 => x"00", -- $0d2a2
          53923 => x"00", -- $0d2a3
          53924 => x"00", -- $0d2a4
          53925 => x"00", -- $0d2a5
          53926 => x"00", -- $0d2a6
          53927 => x"00", -- $0d2a7
          53928 => x"00", -- $0d2a8
          53929 => x"00", -- $0d2a9
          53930 => x"00", -- $0d2aa
          53931 => x"00", -- $0d2ab
          53932 => x"00", -- $0d2ac
          53933 => x"00", -- $0d2ad
          53934 => x"00", -- $0d2ae
          53935 => x"00", -- $0d2af
          53936 => x"00", -- $0d2b0
          53937 => x"00", -- $0d2b1
          53938 => x"00", -- $0d2b2
          53939 => x"00", -- $0d2b3
          53940 => x"00", -- $0d2b4
          53941 => x"00", -- $0d2b5
          53942 => x"00", -- $0d2b6
          53943 => x"00", -- $0d2b7
          53944 => x"00", -- $0d2b8
          53945 => x"00", -- $0d2b9
          53946 => x"00", -- $0d2ba
          53947 => x"00", -- $0d2bb
          53948 => x"00", -- $0d2bc
          53949 => x"00", -- $0d2bd
          53950 => x"00", -- $0d2be
          53951 => x"00", -- $0d2bf
          53952 => x"00", -- $0d2c0
          53953 => x"00", -- $0d2c1
          53954 => x"00", -- $0d2c2
          53955 => x"00", -- $0d2c3
          53956 => x"00", -- $0d2c4
          53957 => x"00", -- $0d2c5
          53958 => x"00", -- $0d2c6
          53959 => x"00", -- $0d2c7
          53960 => x"00", -- $0d2c8
          53961 => x"00", -- $0d2c9
          53962 => x"00", -- $0d2ca
          53963 => x"00", -- $0d2cb
          53964 => x"00", -- $0d2cc
          53965 => x"00", -- $0d2cd
          53966 => x"00", -- $0d2ce
          53967 => x"00", -- $0d2cf
          53968 => x"00", -- $0d2d0
          53969 => x"00", -- $0d2d1
          53970 => x"00", -- $0d2d2
          53971 => x"00", -- $0d2d3
          53972 => x"00", -- $0d2d4
          53973 => x"00", -- $0d2d5
          53974 => x"00", -- $0d2d6
          53975 => x"00", -- $0d2d7
          53976 => x"00", -- $0d2d8
          53977 => x"00", -- $0d2d9
          53978 => x"00", -- $0d2da
          53979 => x"00", -- $0d2db
          53980 => x"00", -- $0d2dc
          53981 => x"00", -- $0d2dd
          53982 => x"00", -- $0d2de
          53983 => x"00", -- $0d2df
          53984 => x"00", -- $0d2e0
          53985 => x"00", -- $0d2e1
          53986 => x"00", -- $0d2e2
          53987 => x"00", -- $0d2e3
          53988 => x"00", -- $0d2e4
          53989 => x"00", -- $0d2e5
          53990 => x"00", -- $0d2e6
          53991 => x"00", -- $0d2e7
          53992 => x"00", -- $0d2e8
          53993 => x"00", -- $0d2e9
          53994 => x"00", -- $0d2ea
          53995 => x"00", -- $0d2eb
          53996 => x"00", -- $0d2ec
          53997 => x"00", -- $0d2ed
          53998 => x"00", -- $0d2ee
          53999 => x"00", -- $0d2ef
          54000 => x"00", -- $0d2f0
          54001 => x"00", -- $0d2f1
          54002 => x"00", -- $0d2f2
          54003 => x"00", -- $0d2f3
          54004 => x"00", -- $0d2f4
          54005 => x"00", -- $0d2f5
          54006 => x"00", -- $0d2f6
          54007 => x"00", -- $0d2f7
          54008 => x"00", -- $0d2f8
          54009 => x"00", -- $0d2f9
          54010 => x"00", -- $0d2fa
          54011 => x"00", -- $0d2fb
          54012 => x"00", -- $0d2fc
          54013 => x"00", -- $0d2fd
          54014 => x"00", -- $0d2fe
          54015 => x"00", -- $0d2ff
          54016 => x"00", -- $0d300
          54017 => x"00", -- $0d301
          54018 => x"00", -- $0d302
          54019 => x"00", -- $0d303
          54020 => x"00", -- $0d304
          54021 => x"00", -- $0d305
          54022 => x"00", -- $0d306
          54023 => x"00", -- $0d307
          54024 => x"00", -- $0d308
          54025 => x"00", -- $0d309
          54026 => x"00", -- $0d30a
          54027 => x"00", -- $0d30b
          54028 => x"00", -- $0d30c
          54029 => x"00", -- $0d30d
          54030 => x"00", -- $0d30e
          54031 => x"00", -- $0d30f
          54032 => x"00", -- $0d310
          54033 => x"00", -- $0d311
          54034 => x"00", -- $0d312
          54035 => x"00", -- $0d313
          54036 => x"00", -- $0d314
          54037 => x"00", -- $0d315
          54038 => x"00", -- $0d316
          54039 => x"00", -- $0d317
          54040 => x"00", -- $0d318
          54041 => x"00", -- $0d319
          54042 => x"00", -- $0d31a
          54043 => x"00", -- $0d31b
          54044 => x"00", -- $0d31c
          54045 => x"00", -- $0d31d
          54046 => x"00", -- $0d31e
          54047 => x"00", -- $0d31f
          54048 => x"00", -- $0d320
          54049 => x"00", -- $0d321
          54050 => x"00", -- $0d322
          54051 => x"00", -- $0d323
          54052 => x"00", -- $0d324
          54053 => x"00", -- $0d325
          54054 => x"00", -- $0d326
          54055 => x"00", -- $0d327
          54056 => x"00", -- $0d328
          54057 => x"00", -- $0d329
          54058 => x"00", -- $0d32a
          54059 => x"00", -- $0d32b
          54060 => x"00", -- $0d32c
          54061 => x"00", -- $0d32d
          54062 => x"00", -- $0d32e
          54063 => x"00", -- $0d32f
          54064 => x"00", -- $0d330
          54065 => x"00", -- $0d331
          54066 => x"00", -- $0d332
          54067 => x"00", -- $0d333
          54068 => x"00", -- $0d334
          54069 => x"00", -- $0d335
          54070 => x"00", -- $0d336
          54071 => x"00", -- $0d337
          54072 => x"00", -- $0d338
          54073 => x"00", -- $0d339
          54074 => x"00", -- $0d33a
          54075 => x"00", -- $0d33b
          54076 => x"00", -- $0d33c
          54077 => x"00", -- $0d33d
          54078 => x"00", -- $0d33e
          54079 => x"00", -- $0d33f
          54080 => x"00", -- $0d340
          54081 => x"00", -- $0d341
          54082 => x"00", -- $0d342
          54083 => x"00", -- $0d343
          54084 => x"00", -- $0d344
          54085 => x"00", -- $0d345
          54086 => x"00", -- $0d346
          54087 => x"00", -- $0d347
          54088 => x"00", -- $0d348
          54089 => x"00", -- $0d349
          54090 => x"00", -- $0d34a
          54091 => x"00", -- $0d34b
          54092 => x"00", -- $0d34c
          54093 => x"00", -- $0d34d
          54094 => x"00", -- $0d34e
          54095 => x"00", -- $0d34f
          54096 => x"00", -- $0d350
          54097 => x"00", -- $0d351
          54098 => x"00", -- $0d352
          54099 => x"00", -- $0d353
          54100 => x"00", -- $0d354
          54101 => x"00", -- $0d355
          54102 => x"00", -- $0d356
          54103 => x"00", -- $0d357
          54104 => x"00", -- $0d358
          54105 => x"00", -- $0d359
          54106 => x"00", -- $0d35a
          54107 => x"00", -- $0d35b
          54108 => x"00", -- $0d35c
          54109 => x"00", -- $0d35d
          54110 => x"00", -- $0d35e
          54111 => x"00", -- $0d35f
          54112 => x"00", -- $0d360
          54113 => x"00", -- $0d361
          54114 => x"00", -- $0d362
          54115 => x"00", -- $0d363
          54116 => x"00", -- $0d364
          54117 => x"00", -- $0d365
          54118 => x"00", -- $0d366
          54119 => x"00", -- $0d367
          54120 => x"00", -- $0d368
          54121 => x"00", -- $0d369
          54122 => x"00", -- $0d36a
          54123 => x"00", -- $0d36b
          54124 => x"00", -- $0d36c
          54125 => x"00", -- $0d36d
          54126 => x"00", -- $0d36e
          54127 => x"00", -- $0d36f
          54128 => x"00", -- $0d370
          54129 => x"00", -- $0d371
          54130 => x"00", -- $0d372
          54131 => x"00", -- $0d373
          54132 => x"00", -- $0d374
          54133 => x"00", -- $0d375
          54134 => x"00", -- $0d376
          54135 => x"00", -- $0d377
          54136 => x"00", -- $0d378
          54137 => x"00", -- $0d379
          54138 => x"00", -- $0d37a
          54139 => x"00", -- $0d37b
          54140 => x"00", -- $0d37c
          54141 => x"00", -- $0d37d
          54142 => x"00", -- $0d37e
          54143 => x"00", -- $0d37f
          54144 => x"00", -- $0d380
          54145 => x"00", -- $0d381
          54146 => x"00", -- $0d382
          54147 => x"00", -- $0d383
          54148 => x"00", -- $0d384
          54149 => x"00", -- $0d385
          54150 => x"00", -- $0d386
          54151 => x"00", -- $0d387
          54152 => x"00", -- $0d388
          54153 => x"00", -- $0d389
          54154 => x"00", -- $0d38a
          54155 => x"00", -- $0d38b
          54156 => x"00", -- $0d38c
          54157 => x"00", -- $0d38d
          54158 => x"00", -- $0d38e
          54159 => x"00", -- $0d38f
          54160 => x"00", -- $0d390
          54161 => x"00", -- $0d391
          54162 => x"00", -- $0d392
          54163 => x"00", -- $0d393
          54164 => x"00", -- $0d394
          54165 => x"00", -- $0d395
          54166 => x"00", -- $0d396
          54167 => x"00", -- $0d397
          54168 => x"00", -- $0d398
          54169 => x"00", -- $0d399
          54170 => x"00", -- $0d39a
          54171 => x"00", -- $0d39b
          54172 => x"00", -- $0d39c
          54173 => x"00", -- $0d39d
          54174 => x"00", -- $0d39e
          54175 => x"00", -- $0d39f
          54176 => x"00", -- $0d3a0
          54177 => x"00", -- $0d3a1
          54178 => x"00", -- $0d3a2
          54179 => x"00", -- $0d3a3
          54180 => x"00", -- $0d3a4
          54181 => x"00", -- $0d3a5
          54182 => x"00", -- $0d3a6
          54183 => x"00", -- $0d3a7
          54184 => x"00", -- $0d3a8
          54185 => x"00", -- $0d3a9
          54186 => x"00", -- $0d3aa
          54187 => x"00", -- $0d3ab
          54188 => x"00", -- $0d3ac
          54189 => x"00", -- $0d3ad
          54190 => x"00", -- $0d3ae
          54191 => x"00", -- $0d3af
          54192 => x"00", -- $0d3b0
          54193 => x"00", -- $0d3b1
          54194 => x"00", -- $0d3b2
          54195 => x"00", -- $0d3b3
          54196 => x"00", -- $0d3b4
          54197 => x"00", -- $0d3b5
          54198 => x"00", -- $0d3b6
          54199 => x"00", -- $0d3b7
          54200 => x"00", -- $0d3b8
          54201 => x"00", -- $0d3b9
          54202 => x"00", -- $0d3ba
          54203 => x"00", -- $0d3bb
          54204 => x"00", -- $0d3bc
          54205 => x"00", -- $0d3bd
          54206 => x"00", -- $0d3be
          54207 => x"00", -- $0d3bf
          54208 => x"00", -- $0d3c0
          54209 => x"00", -- $0d3c1
          54210 => x"00", -- $0d3c2
          54211 => x"00", -- $0d3c3
          54212 => x"00", -- $0d3c4
          54213 => x"00", -- $0d3c5
          54214 => x"00", -- $0d3c6
          54215 => x"00", -- $0d3c7
          54216 => x"00", -- $0d3c8
          54217 => x"00", -- $0d3c9
          54218 => x"00", -- $0d3ca
          54219 => x"00", -- $0d3cb
          54220 => x"00", -- $0d3cc
          54221 => x"00", -- $0d3cd
          54222 => x"00", -- $0d3ce
          54223 => x"00", -- $0d3cf
          54224 => x"00", -- $0d3d0
          54225 => x"00", -- $0d3d1
          54226 => x"00", -- $0d3d2
          54227 => x"00", -- $0d3d3
          54228 => x"00", -- $0d3d4
          54229 => x"00", -- $0d3d5
          54230 => x"00", -- $0d3d6
          54231 => x"00", -- $0d3d7
          54232 => x"00", -- $0d3d8
          54233 => x"00", -- $0d3d9
          54234 => x"00", -- $0d3da
          54235 => x"00", -- $0d3db
          54236 => x"00", -- $0d3dc
          54237 => x"00", -- $0d3dd
          54238 => x"00", -- $0d3de
          54239 => x"00", -- $0d3df
          54240 => x"00", -- $0d3e0
          54241 => x"00", -- $0d3e1
          54242 => x"00", -- $0d3e2
          54243 => x"00", -- $0d3e3
          54244 => x"00", -- $0d3e4
          54245 => x"00", -- $0d3e5
          54246 => x"00", -- $0d3e6
          54247 => x"00", -- $0d3e7
          54248 => x"00", -- $0d3e8
          54249 => x"00", -- $0d3e9
          54250 => x"00", -- $0d3ea
          54251 => x"00", -- $0d3eb
          54252 => x"00", -- $0d3ec
          54253 => x"00", -- $0d3ed
          54254 => x"00", -- $0d3ee
          54255 => x"00", -- $0d3ef
          54256 => x"00", -- $0d3f0
          54257 => x"00", -- $0d3f1
          54258 => x"00", -- $0d3f2
          54259 => x"00", -- $0d3f3
          54260 => x"00", -- $0d3f4
          54261 => x"00", -- $0d3f5
          54262 => x"00", -- $0d3f6
          54263 => x"00", -- $0d3f7
          54264 => x"00", -- $0d3f8
          54265 => x"00", -- $0d3f9
          54266 => x"00", -- $0d3fa
          54267 => x"00", -- $0d3fb
          54268 => x"00", -- $0d3fc
          54269 => x"00", -- $0d3fd
          54270 => x"00", -- $0d3fe
          54271 => x"00", -- $0d3ff
          54272 => x"00", -- $0d400
          54273 => x"00", -- $0d401
          54274 => x"00", -- $0d402
          54275 => x"00", -- $0d403
          54276 => x"00", -- $0d404
          54277 => x"00", -- $0d405
          54278 => x"00", -- $0d406
          54279 => x"00", -- $0d407
          54280 => x"00", -- $0d408
          54281 => x"00", -- $0d409
          54282 => x"00", -- $0d40a
          54283 => x"00", -- $0d40b
          54284 => x"00", -- $0d40c
          54285 => x"00", -- $0d40d
          54286 => x"00", -- $0d40e
          54287 => x"00", -- $0d40f
          54288 => x"00", -- $0d410
          54289 => x"00", -- $0d411
          54290 => x"00", -- $0d412
          54291 => x"00", -- $0d413
          54292 => x"00", -- $0d414
          54293 => x"00", -- $0d415
          54294 => x"00", -- $0d416
          54295 => x"00", -- $0d417
          54296 => x"00", -- $0d418
          54297 => x"00", -- $0d419
          54298 => x"00", -- $0d41a
          54299 => x"00", -- $0d41b
          54300 => x"00", -- $0d41c
          54301 => x"00", -- $0d41d
          54302 => x"00", -- $0d41e
          54303 => x"00", -- $0d41f
          54304 => x"00", -- $0d420
          54305 => x"00", -- $0d421
          54306 => x"00", -- $0d422
          54307 => x"00", -- $0d423
          54308 => x"00", -- $0d424
          54309 => x"00", -- $0d425
          54310 => x"00", -- $0d426
          54311 => x"00", -- $0d427
          54312 => x"00", -- $0d428
          54313 => x"00", -- $0d429
          54314 => x"00", -- $0d42a
          54315 => x"00", -- $0d42b
          54316 => x"00", -- $0d42c
          54317 => x"00", -- $0d42d
          54318 => x"00", -- $0d42e
          54319 => x"00", -- $0d42f
          54320 => x"00", -- $0d430
          54321 => x"00", -- $0d431
          54322 => x"00", -- $0d432
          54323 => x"00", -- $0d433
          54324 => x"00", -- $0d434
          54325 => x"00", -- $0d435
          54326 => x"00", -- $0d436
          54327 => x"00", -- $0d437
          54328 => x"00", -- $0d438
          54329 => x"00", -- $0d439
          54330 => x"00", -- $0d43a
          54331 => x"00", -- $0d43b
          54332 => x"00", -- $0d43c
          54333 => x"00", -- $0d43d
          54334 => x"00", -- $0d43e
          54335 => x"00", -- $0d43f
          54336 => x"00", -- $0d440
          54337 => x"00", -- $0d441
          54338 => x"00", -- $0d442
          54339 => x"00", -- $0d443
          54340 => x"00", -- $0d444
          54341 => x"00", -- $0d445
          54342 => x"00", -- $0d446
          54343 => x"00", -- $0d447
          54344 => x"00", -- $0d448
          54345 => x"00", -- $0d449
          54346 => x"00", -- $0d44a
          54347 => x"00", -- $0d44b
          54348 => x"00", -- $0d44c
          54349 => x"00", -- $0d44d
          54350 => x"00", -- $0d44e
          54351 => x"00", -- $0d44f
          54352 => x"00", -- $0d450
          54353 => x"00", -- $0d451
          54354 => x"00", -- $0d452
          54355 => x"00", -- $0d453
          54356 => x"00", -- $0d454
          54357 => x"00", -- $0d455
          54358 => x"00", -- $0d456
          54359 => x"00", -- $0d457
          54360 => x"00", -- $0d458
          54361 => x"00", -- $0d459
          54362 => x"00", -- $0d45a
          54363 => x"00", -- $0d45b
          54364 => x"00", -- $0d45c
          54365 => x"00", -- $0d45d
          54366 => x"00", -- $0d45e
          54367 => x"00", -- $0d45f
          54368 => x"00", -- $0d460
          54369 => x"00", -- $0d461
          54370 => x"00", -- $0d462
          54371 => x"00", -- $0d463
          54372 => x"00", -- $0d464
          54373 => x"00", -- $0d465
          54374 => x"00", -- $0d466
          54375 => x"00", -- $0d467
          54376 => x"00", -- $0d468
          54377 => x"00", -- $0d469
          54378 => x"00", -- $0d46a
          54379 => x"00", -- $0d46b
          54380 => x"00", -- $0d46c
          54381 => x"00", -- $0d46d
          54382 => x"00", -- $0d46e
          54383 => x"00", -- $0d46f
          54384 => x"00", -- $0d470
          54385 => x"00", -- $0d471
          54386 => x"00", -- $0d472
          54387 => x"00", -- $0d473
          54388 => x"00", -- $0d474
          54389 => x"00", -- $0d475
          54390 => x"00", -- $0d476
          54391 => x"00", -- $0d477
          54392 => x"00", -- $0d478
          54393 => x"00", -- $0d479
          54394 => x"00", -- $0d47a
          54395 => x"00", -- $0d47b
          54396 => x"00", -- $0d47c
          54397 => x"00", -- $0d47d
          54398 => x"00", -- $0d47e
          54399 => x"00", -- $0d47f
          54400 => x"00", -- $0d480
          54401 => x"00", -- $0d481
          54402 => x"00", -- $0d482
          54403 => x"00", -- $0d483
          54404 => x"00", -- $0d484
          54405 => x"00", -- $0d485
          54406 => x"00", -- $0d486
          54407 => x"00", -- $0d487
          54408 => x"00", -- $0d488
          54409 => x"00", -- $0d489
          54410 => x"00", -- $0d48a
          54411 => x"00", -- $0d48b
          54412 => x"00", -- $0d48c
          54413 => x"00", -- $0d48d
          54414 => x"00", -- $0d48e
          54415 => x"00", -- $0d48f
          54416 => x"00", -- $0d490
          54417 => x"00", -- $0d491
          54418 => x"00", -- $0d492
          54419 => x"00", -- $0d493
          54420 => x"00", -- $0d494
          54421 => x"00", -- $0d495
          54422 => x"00", -- $0d496
          54423 => x"00", -- $0d497
          54424 => x"00", -- $0d498
          54425 => x"00", -- $0d499
          54426 => x"00", -- $0d49a
          54427 => x"00", -- $0d49b
          54428 => x"00", -- $0d49c
          54429 => x"00", -- $0d49d
          54430 => x"00", -- $0d49e
          54431 => x"00", -- $0d49f
          54432 => x"00", -- $0d4a0
          54433 => x"00", -- $0d4a1
          54434 => x"00", -- $0d4a2
          54435 => x"00", -- $0d4a3
          54436 => x"00", -- $0d4a4
          54437 => x"00", -- $0d4a5
          54438 => x"00", -- $0d4a6
          54439 => x"00", -- $0d4a7
          54440 => x"00", -- $0d4a8
          54441 => x"00", -- $0d4a9
          54442 => x"00", -- $0d4aa
          54443 => x"00", -- $0d4ab
          54444 => x"00", -- $0d4ac
          54445 => x"00", -- $0d4ad
          54446 => x"00", -- $0d4ae
          54447 => x"00", -- $0d4af
          54448 => x"00", -- $0d4b0
          54449 => x"00", -- $0d4b1
          54450 => x"00", -- $0d4b2
          54451 => x"00", -- $0d4b3
          54452 => x"00", -- $0d4b4
          54453 => x"00", -- $0d4b5
          54454 => x"00", -- $0d4b6
          54455 => x"00", -- $0d4b7
          54456 => x"00", -- $0d4b8
          54457 => x"00", -- $0d4b9
          54458 => x"00", -- $0d4ba
          54459 => x"00", -- $0d4bb
          54460 => x"00", -- $0d4bc
          54461 => x"00", -- $0d4bd
          54462 => x"00", -- $0d4be
          54463 => x"00", -- $0d4bf
          54464 => x"00", -- $0d4c0
          54465 => x"00", -- $0d4c1
          54466 => x"00", -- $0d4c2
          54467 => x"00", -- $0d4c3
          54468 => x"00", -- $0d4c4
          54469 => x"00", -- $0d4c5
          54470 => x"00", -- $0d4c6
          54471 => x"00", -- $0d4c7
          54472 => x"00", -- $0d4c8
          54473 => x"00", -- $0d4c9
          54474 => x"00", -- $0d4ca
          54475 => x"00", -- $0d4cb
          54476 => x"00", -- $0d4cc
          54477 => x"00", -- $0d4cd
          54478 => x"00", -- $0d4ce
          54479 => x"00", -- $0d4cf
          54480 => x"00", -- $0d4d0
          54481 => x"00", -- $0d4d1
          54482 => x"00", -- $0d4d2
          54483 => x"00", -- $0d4d3
          54484 => x"00", -- $0d4d4
          54485 => x"00", -- $0d4d5
          54486 => x"00", -- $0d4d6
          54487 => x"00", -- $0d4d7
          54488 => x"00", -- $0d4d8
          54489 => x"00", -- $0d4d9
          54490 => x"00", -- $0d4da
          54491 => x"00", -- $0d4db
          54492 => x"00", -- $0d4dc
          54493 => x"00", -- $0d4dd
          54494 => x"00", -- $0d4de
          54495 => x"00", -- $0d4df
          54496 => x"00", -- $0d4e0
          54497 => x"00", -- $0d4e1
          54498 => x"00", -- $0d4e2
          54499 => x"00", -- $0d4e3
          54500 => x"00", -- $0d4e4
          54501 => x"00", -- $0d4e5
          54502 => x"00", -- $0d4e6
          54503 => x"00", -- $0d4e7
          54504 => x"00", -- $0d4e8
          54505 => x"00", -- $0d4e9
          54506 => x"00", -- $0d4ea
          54507 => x"00", -- $0d4eb
          54508 => x"00", -- $0d4ec
          54509 => x"00", -- $0d4ed
          54510 => x"00", -- $0d4ee
          54511 => x"00", -- $0d4ef
          54512 => x"00", -- $0d4f0
          54513 => x"00", -- $0d4f1
          54514 => x"00", -- $0d4f2
          54515 => x"00", -- $0d4f3
          54516 => x"00", -- $0d4f4
          54517 => x"00", -- $0d4f5
          54518 => x"00", -- $0d4f6
          54519 => x"00", -- $0d4f7
          54520 => x"00", -- $0d4f8
          54521 => x"00", -- $0d4f9
          54522 => x"00", -- $0d4fa
          54523 => x"00", -- $0d4fb
          54524 => x"00", -- $0d4fc
          54525 => x"00", -- $0d4fd
          54526 => x"00", -- $0d4fe
          54527 => x"00", -- $0d4ff
          54528 => x"00", -- $0d500
          54529 => x"00", -- $0d501
          54530 => x"00", -- $0d502
          54531 => x"00", -- $0d503
          54532 => x"00", -- $0d504
          54533 => x"00", -- $0d505
          54534 => x"00", -- $0d506
          54535 => x"00", -- $0d507
          54536 => x"00", -- $0d508
          54537 => x"00", -- $0d509
          54538 => x"00", -- $0d50a
          54539 => x"00", -- $0d50b
          54540 => x"00", -- $0d50c
          54541 => x"00", -- $0d50d
          54542 => x"00", -- $0d50e
          54543 => x"00", -- $0d50f
          54544 => x"00", -- $0d510
          54545 => x"00", -- $0d511
          54546 => x"00", -- $0d512
          54547 => x"00", -- $0d513
          54548 => x"00", -- $0d514
          54549 => x"00", -- $0d515
          54550 => x"00", -- $0d516
          54551 => x"00", -- $0d517
          54552 => x"00", -- $0d518
          54553 => x"00", -- $0d519
          54554 => x"00", -- $0d51a
          54555 => x"00", -- $0d51b
          54556 => x"00", -- $0d51c
          54557 => x"00", -- $0d51d
          54558 => x"00", -- $0d51e
          54559 => x"00", -- $0d51f
          54560 => x"00", -- $0d520
          54561 => x"00", -- $0d521
          54562 => x"00", -- $0d522
          54563 => x"00", -- $0d523
          54564 => x"00", -- $0d524
          54565 => x"00", -- $0d525
          54566 => x"00", -- $0d526
          54567 => x"00", -- $0d527
          54568 => x"00", -- $0d528
          54569 => x"00", -- $0d529
          54570 => x"00", -- $0d52a
          54571 => x"00", -- $0d52b
          54572 => x"00", -- $0d52c
          54573 => x"00", -- $0d52d
          54574 => x"00", -- $0d52e
          54575 => x"00", -- $0d52f
          54576 => x"00", -- $0d530
          54577 => x"00", -- $0d531
          54578 => x"00", -- $0d532
          54579 => x"00", -- $0d533
          54580 => x"00", -- $0d534
          54581 => x"00", -- $0d535
          54582 => x"00", -- $0d536
          54583 => x"00", -- $0d537
          54584 => x"00", -- $0d538
          54585 => x"00", -- $0d539
          54586 => x"00", -- $0d53a
          54587 => x"00", -- $0d53b
          54588 => x"00", -- $0d53c
          54589 => x"00", -- $0d53d
          54590 => x"00", -- $0d53e
          54591 => x"00", -- $0d53f
          54592 => x"00", -- $0d540
          54593 => x"00", -- $0d541
          54594 => x"00", -- $0d542
          54595 => x"00", -- $0d543
          54596 => x"00", -- $0d544
          54597 => x"00", -- $0d545
          54598 => x"00", -- $0d546
          54599 => x"00", -- $0d547
          54600 => x"00", -- $0d548
          54601 => x"00", -- $0d549
          54602 => x"00", -- $0d54a
          54603 => x"00", -- $0d54b
          54604 => x"00", -- $0d54c
          54605 => x"00", -- $0d54d
          54606 => x"00", -- $0d54e
          54607 => x"00", -- $0d54f
          54608 => x"00", -- $0d550
          54609 => x"00", -- $0d551
          54610 => x"00", -- $0d552
          54611 => x"00", -- $0d553
          54612 => x"00", -- $0d554
          54613 => x"00", -- $0d555
          54614 => x"00", -- $0d556
          54615 => x"00", -- $0d557
          54616 => x"00", -- $0d558
          54617 => x"00", -- $0d559
          54618 => x"00", -- $0d55a
          54619 => x"00", -- $0d55b
          54620 => x"00", -- $0d55c
          54621 => x"00", -- $0d55d
          54622 => x"00", -- $0d55e
          54623 => x"00", -- $0d55f
          54624 => x"00", -- $0d560
          54625 => x"00", -- $0d561
          54626 => x"00", -- $0d562
          54627 => x"00", -- $0d563
          54628 => x"00", -- $0d564
          54629 => x"00", -- $0d565
          54630 => x"00", -- $0d566
          54631 => x"00", -- $0d567
          54632 => x"00", -- $0d568
          54633 => x"00", -- $0d569
          54634 => x"00", -- $0d56a
          54635 => x"00", -- $0d56b
          54636 => x"00", -- $0d56c
          54637 => x"00", -- $0d56d
          54638 => x"00", -- $0d56e
          54639 => x"00", -- $0d56f
          54640 => x"00", -- $0d570
          54641 => x"00", -- $0d571
          54642 => x"00", -- $0d572
          54643 => x"00", -- $0d573
          54644 => x"00", -- $0d574
          54645 => x"00", -- $0d575
          54646 => x"00", -- $0d576
          54647 => x"00", -- $0d577
          54648 => x"00", -- $0d578
          54649 => x"00", -- $0d579
          54650 => x"00", -- $0d57a
          54651 => x"00", -- $0d57b
          54652 => x"00", -- $0d57c
          54653 => x"00", -- $0d57d
          54654 => x"00", -- $0d57e
          54655 => x"00", -- $0d57f
          54656 => x"00", -- $0d580
          54657 => x"00", -- $0d581
          54658 => x"00", -- $0d582
          54659 => x"00", -- $0d583
          54660 => x"00", -- $0d584
          54661 => x"00", -- $0d585
          54662 => x"00", -- $0d586
          54663 => x"00", -- $0d587
          54664 => x"00", -- $0d588
          54665 => x"00", -- $0d589
          54666 => x"00", -- $0d58a
          54667 => x"00", -- $0d58b
          54668 => x"00", -- $0d58c
          54669 => x"00", -- $0d58d
          54670 => x"00", -- $0d58e
          54671 => x"00", -- $0d58f
          54672 => x"00", -- $0d590
          54673 => x"00", -- $0d591
          54674 => x"00", -- $0d592
          54675 => x"00", -- $0d593
          54676 => x"00", -- $0d594
          54677 => x"00", -- $0d595
          54678 => x"00", -- $0d596
          54679 => x"00", -- $0d597
          54680 => x"00", -- $0d598
          54681 => x"00", -- $0d599
          54682 => x"00", -- $0d59a
          54683 => x"00", -- $0d59b
          54684 => x"00", -- $0d59c
          54685 => x"00", -- $0d59d
          54686 => x"00", -- $0d59e
          54687 => x"00", -- $0d59f
          54688 => x"00", -- $0d5a0
          54689 => x"00", -- $0d5a1
          54690 => x"00", -- $0d5a2
          54691 => x"00", -- $0d5a3
          54692 => x"00", -- $0d5a4
          54693 => x"00", -- $0d5a5
          54694 => x"00", -- $0d5a6
          54695 => x"00", -- $0d5a7
          54696 => x"00", -- $0d5a8
          54697 => x"00", -- $0d5a9
          54698 => x"00", -- $0d5aa
          54699 => x"00", -- $0d5ab
          54700 => x"00", -- $0d5ac
          54701 => x"00", -- $0d5ad
          54702 => x"00", -- $0d5ae
          54703 => x"00", -- $0d5af
          54704 => x"00", -- $0d5b0
          54705 => x"00", -- $0d5b1
          54706 => x"00", -- $0d5b2
          54707 => x"00", -- $0d5b3
          54708 => x"00", -- $0d5b4
          54709 => x"00", -- $0d5b5
          54710 => x"00", -- $0d5b6
          54711 => x"00", -- $0d5b7
          54712 => x"00", -- $0d5b8
          54713 => x"00", -- $0d5b9
          54714 => x"00", -- $0d5ba
          54715 => x"00", -- $0d5bb
          54716 => x"00", -- $0d5bc
          54717 => x"00", -- $0d5bd
          54718 => x"00", -- $0d5be
          54719 => x"00", -- $0d5bf
          54720 => x"00", -- $0d5c0
          54721 => x"00", -- $0d5c1
          54722 => x"00", -- $0d5c2
          54723 => x"00", -- $0d5c3
          54724 => x"00", -- $0d5c4
          54725 => x"00", -- $0d5c5
          54726 => x"00", -- $0d5c6
          54727 => x"00", -- $0d5c7
          54728 => x"00", -- $0d5c8
          54729 => x"00", -- $0d5c9
          54730 => x"00", -- $0d5ca
          54731 => x"00", -- $0d5cb
          54732 => x"00", -- $0d5cc
          54733 => x"00", -- $0d5cd
          54734 => x"00", -- $0d5ce
          54735 => x"00", -- $0d5cf
          54736 => x"00", -- $0d5d0
          54737 => x"00", -- $0d5d1
          54738 => x"00", -- $0d5d2
          54739 => x"00", -- $0d5d3
          54740 => x"00", -- $0d5d4
          54741 => x"00", -- $0d5d5
          54742 => x"00", -- $0d5d6
          54743 => x"00", -- $0d5d7
          54744 => x"00", -- $0d5d8
          54745 => x"00", -- $0d5d9
          54746 => x"00", -- $0d5da
          54747 => x"00", -- $0d5db
          54748 => x"00", -- $0d5dc
          54749 => x"00", -- $0d5dd
          54750 => x"00", -- $0d5de
          54751 => x"00", -- $0d5df
          54752 => x"00", -- $0d5e0
          54753 => x"00", -- $0d5e1
          54754 => x"00", -- $0d5e2
          54755 => x"00", -- $0d5e3
          54756 => x"00", -- $0d5e4
          54757 => x"00", -- $0d5e5
          54758 => x"00", -- $0d5e6
          54759 => x"00", -- $0d5e7
          54760 => x"00", -- $0d5e8
          54761 => x"00", -- $0d5e9
          54762 => x"00", -- $0d5ea
          54763 => x"00", -- $0d5eb
          54764 => x"00", -- $0d5ec
          54765 => x"00", -- $0d5ed
          54766 => x"00", -- $0d5ee
          54767 => x"00", -- $0d5ef
          54768 => x"00", -- $0d5f0
          54769 => x"00", -- $0d5f1
          54770 => x"00", -- $0d5f2
          54771 => x"00", -- $0d5f3
          54772 => x"00", -- $0d5f4
          54773 => x"00", -- $0d5f5
          54774 => x"00", -- $0d5f6
          54775 => x"00", -- $0d5f7
          54776 => x"00", -- $0d5f8
          54777 => x"00", -- $0d5f9
          54778 => x"00", -- $0d5fa
          54779 => x"00", -- $0d5fb
          54780 => x"00", -- $0d5fc
          54781 => x"00", -- $0d5fd
          54782 => x"00", -- $0d5fe
          54783 => x"00", -- $0d5ff
          54784 => x"00", -- $0d600
          54785 => x"00", -- $0d601
          54786 => x"00", -- $0d602
          54787 => x"00", -- $0d603
          54788 => x"00", -- $0d604
          54789 => x"00", -- $0d605
          54790 => x"00", -- $0d606
          54791 => x"00", -- $0d607
          54792 => x"00", -- $0d608
          54793 => x"00", -- $0d609
          54794 => x"00", -- $0d60a
          54795 => x"00", -- $0d60b
          54796 => x"00", -- $0d60c
          54797 => x"00", -- $0d60d
          54798 => x"00", -- $0d60e
          54799 => x"00", -- $0d60f
          54800 => x"00", -- $0d610
          54801 => x"00", -- $0d611
          54802 => x"00", -- $0d612
          54803 => x"00", -- $0d613
          54804 => x"00", -- $0d614
          54805 => x"00", -- $0d615
          54806 => x"00", -- $0d616
          54807 => x"00", -- $0d617
          54808 => x"00", -- $0d618
          54809 => x"00", -- $0d619
          54810 => x"00", -- $0d61a
          54811 => x"00", -- $0d61b
          54812 => x"00", -- $0d61c
          54813 => x"00", -- $0d61d
          54814 => x"00", -- $0d61e
          54815 => x"00", -- $0d61f
          54816 => x"00", -- $0d620
          54817 => x"00", -- $0d621
          54818 => x"00", -- $0d622
          54819 => x"00", -- $0d623
          54820 => x"00", -- $0d624
          54821 => x"00", -- $0d625
          54822 => x"00", -- $0d626
          54823 => x"00", -- $0d627
          54824 => x"00", -- $0d628
          54825 => x"00", -- $0d629
          54826 => x"00", -- $0d62a
          54827 => x"00", -- $0d62b
          54828 => x"00", -- $0d62c
          54829 => x"00", -- $0d62d
          54830 => x"00", -- $0d62e
          54831 => x"00", -- $0d62f
          54832 => x"00", -- $0d630
          54833 => x"00", -- $0d631
          54834 => x"00", -- $0d632
          54835 => x"00", -- $0d633
          54836 => x"00", -- $0d634
          54837 => x"00", -- $0d635
          54838 => x"00", -- $0d636
          54839 => x"00", -- $0d637
          54840 => x"00", -- $0d638
          54841 => x"00", -- $0d639
          54842 => x"00", -- $0d63a
          54843 => x"00", -- $0d63b
          54844 => x"00", -- $0d63c
          54845 => x"00", -- $0d63d
          54846 => x"00", -- $0d63e
          54847 => x"00", -- $0d63f
          54848 => x"00", -- $0d640
          54849 => x"00", -- $0d641
          54850 => x"00", -- $0d642
          54851 => x"00", -- $0d643
          54852 => x"00", -- $0d644
          54853 => x"00", -- $0d645
          54854 => x"00", -- $0d646
          54855 => x"00", -- $0d647
          54856 => x"00", -- $0d648
          54857 => x"00", -- $0d649
          54858 => x"00", -- $0d64a
          54859 => x"00", -- $0d64b
          54860 => x"00", -- $0d64c
          54861 => x"00", -- $0d64d
          54862 => x"00", -- $0d64e
          54863 => x"00", -- $0d64f
          54864 => x"00", -- $0d650
          54865 => x"00", -- $0d651
          54866 => x"00", -- $0d652
          54867 => x"00", -- $0d653
          54868 => x"00", -- $0d654
          54869 => x"00", -- $0d655
          54870 => x"00", -- $0d656
          54871 => x"00", -- $0d657
          54872 => x"00", -- $0d658
          54873 => x"00", -- $0d659
          54874 => x"00", -- $0d65a
          54875 => x"00", -- $0d65b
          54876 => x"00", -- $0d65c
          54877 => x"00", -- $0d65d
          54878 => x"00", -- $0d65e
          54879 => x"00", -- $0d65f
          54880 => x"00", -- $0d660
          54881 => x"00", -- $0d661
          54882 => x"00", -- $0d662
          54883 => x"00", -- $0d663
          54884 => x"00", -- $0d664
          54885 => x"00", -- $0d665
          54886 => x"00", -- $0d666
          54887 => x"00", -- $0d667
          54888 => x"00", -- $0d668
          54889 => x"00", -- $0d669
          54890 => x"00", -- $0d66a
          54891 => x"00", -- $0d66b
          54892 => x"00", -- $0d66c
          54893 => x"00", -- $0d66d
          54894 => x"00", -- $0d66e
          54895 => x"00", -- $0d66f
          54896 => x"00", -- $0d670
          54897 => x"00", -- $0d671
          54898 => x"00", -- $0d672
          54899 => x"00", -- $0d673
          54900 => x"00", -- $0d674
          54901 => x"00", -- $0d675
          54902 => x"00", -- $0d676
          54903 => x"00", -- $0d677
          54904 => x"00", -- $0d678
          54905 => x"00", -- $0d679
          54906 => x"00", -- $0d67a
          54907 => x"00", -- $0d67b
          54908 => x"00", -- $0d67c
          54909 => x"00", -- $0d67d
          54910 => x"00", -- $0d67e
          54911 => x"00", -- $0d67f
          54912 => x"00", -- $0d680
          54913 => x"00", -- $0d681
          54914 => x"00", -- $0d682
          54915 => x"00", -- $0d683
          54916 => x"00", -- $0d684
          54917 => x"00", -- $0d685
          54918 => x"00", -- $0d686
          54919 => x"00", -- $0d687
          54920 => x"00", -- $0d688
          54921 => x"00", -- $0d689
          54922 => x"00", -- $0d68a
          54923 => x"00", -- $0d68b
          54924 => x"00", -- $0d68c
          54925 => x"00", -- $0d68d
          54926 => x"00", -- $0d68e
          54927 => x"00", -- $0d68f
          54928 => x"00", -- $0d690
          54929 => x"00", -- $0d691
          54930 => x"00", -- $0d692
          54931 => x"00", -- $0d693
          54932 => x"00", -- $0d694
          54933 => x"00", -- $0d695
          54934 => x"00", -- $0d696
          54935 => x"00", -- $0d697
          54936 => x"00", -- $0d698
          54937 => x"00", -- $0d699
          54938 => x"00", -- $0d69a
          54939 => x"00", -- $0d69b
          54940 => x"00", -- $0d69c
          54941 => x"00", -- $0d69d
          54942 => x"00", -- $0d69e
          54943 => x"00", -- $0d69f
          54944 => x"00", -- $0d6a0
          54945 => x"00", -- $0d6a1
          54946 => x"00", -- $0d6a2
          54947 => x"00", -- $0d6a3
          54948 => x"00", -- $0d6a4
          54949 => x"00", -- $0d6a5
          54950 => x"00", -- $0d6a6
          54951 => x"00", -- $0d6a7
          54952 => x"00", -- $0d6a8
          54953 => x"00", -- $0d6a9
          54954 => x"00", -- $0d6aa
          54955 => x"00", -- $0d6ab
          54956 => x"00", -- $0d6ac
          54957 => x"00", -- $0d6ad
          54958 => x"00", -- $0d6ae
          54959 => x"00", -- $0d6af
          54960 => x"00", -- $0d6b0
          54961 => x"00", -- $0d6b1
          54962 => x"00", -- $0d6b2
          54963 => x"00", -- $0d6b3
          54964 => x"00", -- $0d6b4
          54965 => x"00", -- $0d6b5
          54966 => x"00", -- $0d6b6
          54967 => x"00", -- $0d6b7
          54968 => x"00", -- $0d6b8
          54969 => x"00", -- $0d6b9
          54970 => x"00", -- $0d6ba
          54971 => x"00", -- $0d6bb
          54972 => x"00", -- $0d6bc
          54973 => x"00", -- $0d6bd
          54974 => x"00", -- $0d6be
          54975 => x"00", -- $0d6bf
          54976 => x"00", -- $0d6c0
          54977 => x"00", -- $0d6c1
          54978 => x"00", -- $0d6c2
          54979 => x"00", -- $0d6c3
          54980 => x"00", -- $0d6c4
          54981 => x"00", -- $0d6c5
          54982 => x"00", -- $0d6c6
          54983 => x"00", -- $0d6c7
          54984 => x"00", -- $0d6c8
          54985 => x"00", -- $0d6c9
          54986 => x"00", -- $0d6ca
          54987 => x"00", -- $0d6cb
          54988 => x"00", -- $0d6cc
          54989 => x"00", -- $0d6cd
          54990 => x"00", -- $0d6ce
          54991 => x"00", -- $0d6cf
          54992 => x"00", -- $0d6d0
          54993 => x"00", -- $0d6d1
          54994 => x"00", -- $0d6d2
          54995 => x"00", -- $0d6d3
          54996 => x"00", -- $0d6d4
          54997 => x"00", -- $0d6d5
          54998 => x"00", -- $0d6d6
          54999 => x"00", -- $0d6d7
          55000 => x"00", -- $0d6d8
          55001 => x"00", -- $0d6d9
          55002 => x"00", -- $0d6da
          55003 => x"00", -- $0d6db
          55004 => x"00", -- $0d6dc
          55005 => x"00", -- $0d6dd
          55006 => x"00", -- $0d6de
          55007 => x"00", -- $0d6df
          55008 => x"00", -- $0d6e0
          55009 => x"00", -- $0d6e1
          55010 => x"00", -- $0d6e2
          55011 => x"00", -- $0d6e3
          55012 => x"00", -- $0d6e4
          55013 => x"00", -- $0d6e5
          55014 => x"00", -- $0d6e6
          55015 => x"00", -- $0d6e7
          55016 => x"00", -- $0d6e8
          55017 => x"00", -- $0d6e9
          55018 => x"00", -- $0d6ea
          55019 => x"00", -- $0d6eb
          55020 => x"00", -- $0d6ec
          55021 => x"00", -- $0d6ed
          55022 => x"00", -- $0d6ee
          55023 => x"00", -- $0d6ef
          55024 => x"00", -- $0d6f0
          55025 => x"00", -- $0d6f1
          55026 => x"00", -- $0d6f2
          55027 => x"00", -- $0d6f3
          55028 => x"00", -- $0d6f4
          55029 => x"00", -- $0d6f5
          55030 => x"00", -- $0d6f6
          55031 => x"00", -- $0d6f7
          55032 => x"00", -- $0d6f8
          55033 => x"00", -- $0d6f9
          55034 => x"00", -- $0d6fa
          55035 => x"00", -- $0d6fb
          55036 => x"00", -- $0d6fc
          55037 => x"00", -- $0d6fd
          55038 => x"00", -- $0d6fe
          55039 => x"00", -- $0d6ff
          55040 => x"00", -- $0d700
          55041 => x"00", -- $0d701
          55042 => x"00", -- $0d702
          55043 => x"00", -- $0d703
          55044 => x"00", -- $0d704
          55045 => x"00", -- $0d705
          55046 => x"00", -- $0d706
          55047 => x"00", -- $0d707
          55048 => x"00", -- $0d708
          55049 => x"00", -- $0d709
          55050 => x"00", -- $0d70a
          55051 => x"00", -- $0d70b
          55052 => x"00", -- $0d70c
          55053 => x"00", -- $0d70d
          55054 => x"00", -- $0d70e
          55055 => x"00", -- $0d70f
          55056 => x"00", -- $0d710
          55057 => x"00", -- $0d711
          55058 => x"00", -- $0d712
          55059 => x"00", -- $0d713
          55060 => x"00", -- $0d714
          55061 => x"00", -- $0d715
          55062 => x"00", -- $0d716
          55063 => x"00", -- $0d717
          55064 => x"00", -- $0d718
          55065 => x"00", -- $0d719
          55066 => x"00", -- $0d71a
          55067 => x"00", -- $0d71b
          55068 => x"00", -- $0d71c
          55069 => x"00", -- $0d71d
          55070 => x"00", -- $0d71e
          55071 => x"00", -- $0d71f
          55072 => x"00", -- $0d720
          55073 => x"00", -- $0d721
          55074 => x"00", -- $0d722
          55075 => x"00", -- $0d723
          55076 => x"00", -- $0d724
          55077 => x"00", -- $0d725
          55078 => x"00", -- $0d726
          55079 => x"00", -- $0d727
          55080 => x"00", -- $0d728
          55081 => x"00", -- $0d729
          55082 => x"00", -- $0d72a
          55083 => x"00", -- $0d72b
          55084 => x"00", -- $0d72c
          55085 => x"00", -- $0d72d
          55086 => x"00", -- $0d72e
          55087 => x"00", -- $0d72f
          55088 => x"00", -- $0d730
          55089 => x"00", -- $0d731
          55090 => x"00", -- $0d732
          55091 => x"00", -- $0d733
          55092 => x"00", -- $0d734
          55093 => x"00", -- $0d735
          55094 => x"00", -- $0d736
          55095 => x"00", -- $0d737
          55096 => x"00", -- $0d738
          55097 => x"00", -- $0d739
          55098 => x"00", -- $0d73a
          55099 => x"00", -- $0d73b
          55100 => x"00", -- $0d73c
          55101 => x"00", -- $0d73d
          55102 => x"00", -- $0d73e
          55103 => x"00", -- $0d73f
          55104 => x"00", -- $0d740
          55105 => x"00", -- $0d741
          55106 => x"00", -- $0d742
          55107 => x"00", -- $0d743
          55108 => x"00", -- $0d744
          55109 => x"00", -- $0d745
          55110 => x"00", -- $0d746
          55111 => x"00", -- $0d747
          55112 => x"00", -- $0d748
          55113 => x"00", -- $0d749
          55114 => x"00", -- $0d74a
          55115 => x"00", -- $0d74b
          55116 => x"00", -- $0d74c
          55117 => x"00", -- $0d74d
          55118 => x"00", -- $0d74e
          55119 => x"00", -- $0d74f
          55120 => x"00", -- $0d750
          55121 => x"00", -- $0d751
          55122 => x"00", -- $0d752
          55123 => x"00", -- $0d753
          55124 => x"00", -- $0d754
          55125 => x"00", -- $0d755
          55126 => x"00", -- $0d756
          55127 => x"00", -- $0d757
          55128 => x"00", -- $0d758
          55129 => x"00", -- $0d759
          55130 => x"00", -- $0d75a
          55131 => x"00", -- $0d75b
          55132 => x"00", -- $0d75c
          55133 => x"00", -- $0d75d
          55134 => x"00", -- $0d75e
          55135 => x"00", -- $0d75f
          55136 => x"00", -- $0d760
          55137 => x"00", -- $0d761
          55138 => x"00", -- $0d762
          55139 => x"00", -- $0d763
          55140 => x"00", -- $0d764
          55141 => x"00", -- $0d765
          55142 => x"00", -- $0d766
          55143 => x"00", -- $0d767
          55144 => x"00", -- $0d768
          55145 => x"00", -- $0d769
          55146 => x"00", -- $0d76a
          55147 => x"00", -- $0d76b
          55148 => x"00", -- $0d76c
          55149 => x"00", -- $0d76d
          55150 => x"00", -- $0d76e
          55151 => x"00", -- $0d76f
          55152 => x"00", -- $0d770
          55153 => x"00", -- $0d771
          55154 => x"00", -- $0d772
          55155 => x"00", -- $0d773
          55156 => x"00", -- $0d774
          55157 => x"00", -- $0d775
          55158 => x"00", -- $0d776
          55159 => x"00", -- $0d777
          55160 => x"00", -- $0d778
          55161 => x"00", -- $0d779
          55162 => x"00", -- $0d77a
          55163 => x"00", -- $0d77b
          55164 => x"00", -- $0d77c
          55165 => x"00", -- $0d77d
          55166 => x"00", -- $0d77e
          55167 => x"00", -- $0d77f
          55168 => x"00", -- $0d780
          55169 => x"00", -- $0d781
          55170 => x"00", -- $0d782
          55171 => x"00", -- $0d783
          55172 => x"00", -- $0d784
          55173 => x"00", -- $0d785
          55174 => x"00", -- $0d786
          55175 => x"00", -- $0d787
          55176 => x"00", -- $0d788
          55177 => x"00", -- $0d789
          55178 => x"00", -- $0d78a
          55179 => x"00", -- $0d78b
          55180 => x"00", -- $0d78c
          55181 => x"00", -- $0d78d
          55182 => x"00", -- $0d78e
          55183 => x"00", -- $0d78f
          55184 => x"00", -- $0d790
          55185 => x"00", -- $0d791
          55186 => x"00", -- $0d792
          55187 => x"00", -- $0d793
          55188 => x"00", -- $0d794
          55189 => x"00", -- $0d795
          55190 => x"00", -- $0d796
          55191 => x"00", -- $0d797
          55192 => x"00", -- $0d798
          55193 => x"00", -- $0d799
          55194 => x"00", -- $0d79a
          55195 => x"00", -- $0d79b
          55196 => x"00", -- $0d79c
          55197 => x"00", -- $0d79d
          55198 => x"00", -- $0d79e
          55199 => x"00", -- $0d79f
          55200 => x"00", -- $0d7a0
          55201 => x"00", -- $0d7a1
          55202 => x"00", -- $0d7a2
          55203 => x"00", -- $0d7a3
          55204 => x"00", -- $0d7a4
          55205 => x"00", -- $0d7a5
          55206 => x"00", -- $0d7a6
          55207 => x"00", -- $0d7a7
          55208 => x"00", -- $0d7a8
          55209 => x"00", -- $0d7a9
          55210 => x"00", -- $0d7aa
          55211 => x"00", -- $0d7ab
          55212 => x"00", -- $0d7ac
          55213 => x"00", -- $0d7ad
          55214 => x"00", -- $0d7ae
          55215 => x"00", -- $0d7af
          55216 => x"00", -- $0d7b0
          55217 => x"00", -- $0d7b1
          55218 => x"00", -- $0d7b2
          55219 => x"00", -- $0d7b3
          55220 => x"00", -- $0d7b4
          55221 => x"00", -- $0d7b5
          55222 => x"00", -- $0d7b6
          55223 => x"00", -- $0d7b7
          55224 => x"00", -- $0d7b8
          55225 => x"00", -- $0d7b9
          55226 => x"00", -- $0d7ba
          55227 => x"00", -- $0d7bb
          55228 => x"00", -- $0d7bc
          55229 => x"00", -- $0d7bd
          55230 => x"00", -- $0d7be
          55231 => x"00", -- $0d7bf
          55232 => x"00", -- $0d7c0
          55233 => x"00", -- $0d7c1
          55234 => x"00", -- $0d7c2
          55235 => x"00", -- $0d7c3
          55236 => x"00", -- $0d7c4
          55237 => x"00", -- $0d7c5
          55238 => x"00", -- $0d7c6
          55239 => x"00", -- $0d7c7
          55240 => x"00", -- $0d7c8
          55241 => x"00", -- $0d7c9
          55242 => x"00", -- $0d7ca
          55243 => x"00", -- $0d7cb
          55244 => x"00", -- $0d7cc
          55245 => x"00", -- $0d7cd
          55246 => x"00", -- $0d7ce
          55247 => x"00", -- $0d7cf
          55248 => x"00", -- $0d7d0
          55249 => x"00", -- $0d7d1
          55250 => x"00", -- $0d7d2
          55251 => x"00", -- $0d7d3
          55252 => x"00", -- $0d7d4
          55253 => x"00", -- $0d7d5
          55254 => x"00", -- $0d7d6
          55255 => x"00", -- $0d7d7
          55256 => x"00", -- $0d7d8
          55257 => x"00", -- $0d7d9
          55258 => x"00", -- $0d7da
          55259 => x"00", -- $0d7db
          55260 => x"00", -- $0d7dc
          55261 => x"00", -- $0d7dd
          55262 => x"00", -- $0d7de
          55263 => x"00", -- $0d7df
          55264 => x"00", -- $0d7e0
          55265 => x"00", -- $0d7e1
          55266 => x"00", -- $0d7e2
          55267 => x"00", -- $0d7e3
          55268 => x"00", -- $0d7e4
          55269 => x"00", -- $0d7e5
          55270 => x"00", -- $0d7e6
          55271 => x"00", -- $0d7e7
          55272 => x"00", -- $0d7e8
          55273 => x"00", -- $0d7e9
          55274 => x"00", -- $0d7ea
          55275 => x"00", -- $0d7eb
          55276 => x"00", -- $0d7ec
          55277 => x"00", -- $0d7ed
          55278 => x"00", -- $0d7ee
          55279 => x"00", -- $0d7ef
          55280 => x"00", -- $0d7f0
          55281 => x"00", -- $0d7f1
          55282 => x"00", -- $0d7f2
          55283 => x"00", -- $0d7f3
          55284 => x"00", -- $0d7f4
          55285 => x"00", -- $0d7f5
          55286 => x"00", -- $0d7f6
          55287 => x"00", -- $0d7f7
          55288 => x"00", -- $0d7f8
          55289 => x"00", -- $0d7f9
          55290 => x"00", -- $0d7fa
          55291 => x"00", -- $0d7fb
          55292 => x"00", -- $0d7fc
          55293 => x"00", -- $0d7fd
          55294 => x"00", -- $0d7fe
          55295 => x"00", -- $0d7ff
          55296 => x"00", -- $0d800
          55297 => x"00", -- $0d801
          55298 => x"00", -- $0d802
          55299 => x"00", -- $0d803
          55300 => x"00", -- $0d804
          55301 => x"00", -- $0d805
          55302 => x"00", -- $0d806
          55303 => x"00", -- $0d807
          55304 => x"00", -- $0d808
          55305 => x"00", -- $0d809
          55306 => x"00", -- $0d80a
          55307 => x"00", -- $0d80b
          55308 => x"00", -- $0d80c
          55309 => x"00", -- $0d80d
          55310 => x"00", -- $0d80e
          55311 => x"00", -- $0d80f
          55312 => x"00", -- $0d810
          55313 => x"00", -- $0d811
          55314 => x"00", -- $0d812
          55315 => x"00", -- $0d813
          55316 => x"00", -- $0d814
          55317 => x"00", -- $0d815
          55318 => x"00", -- $0d816
          55319 => x"00", -- $0d817
          55320 => x"00", -- $0d818
          55321 => x"00", -- $0d819
          55322 => x"00", -- $0d81a
          55323 => x"00", -- $0d81b
          55324 => x"00", -- $0d81c
          55325 => x"00", -- $0d81d
          55326 => x"00", -- $0d81e
          55327 => x"00", -- $0d81f
          55328 => x"00", -- $0d820
          55329 => x"00", -- $0d821
          55330 => x"00", -- $0d822
          55331 => x"00", -- $0d823
          55332 => x"00", -- $0d824
          55333 => x"00", -- $0d825
          55334 => x"00", -- $0d826
          55335 => x"00", -- $0d827
          55336 => x"00", -- $0d828
          55337 => x"00", -- $0d829
          55338 => x"00", -- $0d82a
          55339 => x"00", -- $0d82b
          55340 => x"00", -- $0d82c
          55341 => x"00", -- $0d82d
          55342 => x"00", -- $0d82e
          55343 => x"00", -- $0d82f
          55344 => x"00", -- $0d830
          55345 => x"00", -- $0d831
          55346 => x"00", -- $0d832
          55347 => x"00", -- $0d833
          55348 => x"00", -- $0d834
          55349 => x"00", -- $0d835
          55350 => x"00", -- $0d836
          55351 => x"00", -- $0d837
          55352 => x"00", -- $0d838
          55353 => x"00", -- $0d839
          55354 => x"00", -- $0d83a
          55355 => x"00", -- $0d83b
          55356 => x"00", -- $0d83c
          55357 => x"00", -- $0d83d
          55358 => x"00", -- $0d83e
          55359 => x"00", -- $0d83f
          55360 => x"00", -- $0d840
          55361 => x"00", -- $0d841
          55362 => x"00", -- $0d842
          55363 => x"00", -- $0d843
          55364 => x"00", -- $0d844
          55365 => x"00", -- $0d845
          55366 => x"00", -- $0d846
          55367 => x"00", -- $0d847
          55368 => x"00", -- $0d848
          55369 => x"00", -- $0d849
          55370 => x"00", -- $0d84a
          55371 => x"00", -- $0d84b
          55372 => x"00", -- $0d84c
          55373 => x"00", -- $0d84d
          55374 => x"00", -- $0d84e
          55375 => x"00", -- $0d84f
          55376 => x"00", -- $0d850
          55377 => x"00", -- $0d851
          55378 => x"00", -- $0d852
          55379 => x"00", -- $0d853
          55380 => x"00", -- $0d854
          55381 => x"00", -- $0d855
          55382 => x"00", -- $0d856
          55383 => x"00", -- $0d857
          55384 => x"00", -- $0d858
          55385 => x"00", -- $0d859
          55386 => x"00", -- $0d85a
          55387 => x"00", -- $0d85b
          55388 => x"00", -- $0d85c
          55389 => x"00", -- $0d85d
          55390 => x"00", -- $0d85e
          55391 => x"00", -- $0d85f
          55392 => x"00", -- $0d860
          55393 => x"00", -- $0d861
          55394 => x"00", -- $0d862
          55395 => x"00", -- $0d863
          55396 => x"00", -- $0d864
          55397 => x"00", -- $0d865
          55398 => x"00", -- $0d866
          55399 => x"00", -- $0d867
          55400 => x"00", -- $0d868
          55401 => x"00", -- $0d869
          55402 => x"00", -- $0d86a
          55403 => x"00", -- $0d86b
          55404 => x"00", -- $0d86c
          55405 => x"00", -- $0d86d
          55406 => x"00", -- $0d86e
          55407 => x"00", -- $0d86f
          55408 => x"00", -- $0d870
          55409 => x"00", -- $0d871
          55410 => x"00", -- $0d872
          55411 => x"00", -- $0d873
          55412 => x"00", -- $0d874
          55413 => x"00", -- $0d875
          55414 => x"00", -- $0d876
          55415 => x"00", -- $0d877
          55416 => x"00", -- $0d878
          55417 => x"00", -- $0d879
          55418 => x"00", -- $0d87a
          55419 => x"00", -- $0d87b
          55420 => x"00", -- $0d87c
          55421 => x"00", -- $0d87d
          55422 => x"00", -- $0d87e
          55423 => x"00", -- $0d87f
          55424 => x"00", -- $0d880
          55425 => x"00", -- $0d881
          55426 => x"00", -- $0d882
          55427 => x"00", -- $0d883
          55428 => x"00", -- $0d884
          55429 => x"00", -- $0d885
          55430 => x"00", -- $0d886
          55431 => x"00", -- $0d887
          55432 => x"00", -- $0d888
          55433 => x"00", -- $0d889
          55434 => x"00", -- $0d88a
          55435 => x"00", -- $0d88b
          55436 => x"00", -- $0d88c
          55437 => x"00", -- $0d88d
          55438 => x"00", -- $0d88e
          55439 => x"00", -- $0d88f
          55440 => x"00", -- $0d890
          55441 => x"00", -- $0d891
          55442 => x"00", -- $0d892
          55443 => x"00", -- $0d893
          55444 => x"00", -- $0d894
          55445 => x"00", -- $0d895
          55446 => x"00", -- $0d896
          55447 => x"00", -- $0d897
          55448 => x"00", -- $0d898
          55449 => x"00", -- $0d899
          55450 => x"00", -- $0d89a
          55451 => x"00", -- $0d89b
          55452 => x"00", -- $0d89c
          55453 => x"00", -- $0d89d
          55454 => x"00", -- $0d89e
          55455 => x"00", -- $0d89f
          55456 => x"00", -- $0d8a0
          55457 => x"00", -- $0d8a1
          55458 => x"00", -- $0d8a2
          55459 => x"00", -- $0d8a3
          55460 => x"00", -- $0d8a4
          55461 => x"00", -- $0d8a5
          55462 => x"00", -- $0d8a6
          55463 => x"00", -- $0d8a7
          55464 => x"00", -- $0d8a8
          55465 => x"00", -- $0d8a9
          55466 => x"00", -- $0d8aa
          55467 => x"00", -- $0d8ab
          55468 => x"00", -- $0d8ac
          55469 => x"00", -- $0d8ad
          55470 => x"00", -- $0d8ae
          55471 => x"00", -- $0d8af
          55472 => x"00", -- $0d8b0
          55473 => x"00", -- $0d8b1
          55474 => x"00", -- $0d8b2
          55475 => x"00", -- $0d8b3
          55476 => x"00", -- $0d8b4
          55477 => x"00", -- $0d8b5
          55478 => x"00", -- $0d8b6
          55479 => x"00", -- $0d8b7
          55480 => x"00", -- $0d8b8
          55481 => x"00", -- $0d8b9
          55482 => x"00", -- $0d8ba
          55483 => x"00", -- $0d8bb
          55484 => x"00", -- $0d8bc
          55485 => x"00", -- $0d8bd
          55486 => x"00", -- $0d8be
          55487 => x"00", -- $0d8bf
          55488 => x"00", -- $0d8c0
          55489 => x"00", -- $0d8c1
          55490 => x"00", -- $0d8c2
          55491 => x"00", -- $0d8c3
          55492 => x"00", -- $0d8c4
          55493 => x"00", -- $0d8c5
          55494 => x"00", -- $0d8c6
          55495 => x"00", -- $0d8c7
          55496 => x"00", -- $0d8c8
          55497 => x"00", -- $0d8c9
          55498 => x"00", -- $0d8ca
          55499 => x"00", -- $0d8cb
          55500 => x"00", -- $0d8cc
          55501 => x"00", -- $0d8cd
          55502 => x"00", -- $0d8ce
          55503 => x"00", -- $0d8cf
          55504 => x"00", -- $0d8d0
          55505 => x"00", -- $0d8d1
          55506 => x"00", -- $0d8d2
          55507 => x"00", -- $0d8d3
          55508 => x"00", -- $0d8d4
          55509 => x"00", -- $0d8d5
          55510 => x"00", -- $0d8d6
          55511 => x"00", -- $0d8d7
          55512 => x"00", -- $0d8d8
          55513 => x"00", -- $0d8d9
          55514 => x"00", -- $0d8da
          55515 => x"00", -- $0d8db
          55516 => x"00", -- $0d8dc
          55517 => x"00", -- $0d8dd
          55518 => x"00", -- $0d8de
          55519 => x"00", -- $0d8df
          55520 => x"00", -- $0d8e0
          55521 => x"00", -- $0d8e1
          55522 => x"00", -- $0d8e2
          55523 => x"00", -- $0d8e3
          55524 => x"00", -- $0d8e4
          55525 => x"00", -- $0d8e5
          55526 => x"00", -- $0d8e6
          55527 => x"00", -- $0d8e7
          55528 => x"00", -- $0d8e8
          55529 => x"00", -- $0d8e9
          55530 => x"00", -- $0d8ea
          55531 => x"00", -- $0d8eb
          55532 => x"00", -- $0d8ec
          55533 => x"00", -- $0d8ed
          55534 => x"00", -- $0d8ee
          55535 => x"00", -- $0d8ef
          55536 => x"00", -- $0d8f0
          55537 => x"00", -- $0d8f1
          55538 => x"00", -- $0d8f2
          55539 => x"00", -- $0d8f3
          55540 => x"00", -- $0d8f4
          55541 => x"00", -- $0d8f5
          55542 => x"00", -- $0d8f6
          55543 => x"00", -- $0d8f7
          55544 => x"00", -- $0d8f8
          55545 => x"00", -- $0d8f9
          55546 => x"00", -- $0d8fa
          55547 => x"00", -- $0d8fb
          55548 => x"00", -- $0d8fc
          55549 => x"00", -- $0d8fd
          55550 => x"00", -- $0d8fe
          55551 => x"00", -- $0d8ff
          55552 => x"00", -- $0d900
          55553 => x"00", -- $0d901
          55554 => x"00", -- $0d902
          55555 => x"00", -- $0d903
          55556 => x"00", -- $0d904
          55557 => x"00", -- $0d905
          55558 => x"00", -- $0d906
          55559 => x"00", -- $0d907
          55560 => x"00", -- $0d908
          55561 => x"00", -- $0d909
          55562 => x"00", -- $0d90a
          55563 => x"00", -- $0d90b
          55564 => x"00", -- $0d90c
          55565 => x"00", -- $0d90d
          55566 => x"00", -- $0d90e
          55567 => x"00", -- $0d90f
          55568 => x"00", -- $0d910
          55569 => x"00", -- $0d911
          55570 => x"00", -- $0d912
          55571 => x"00", -- $0d913
          55572 => x"00", -- $0d914
          55573 => x"00", -- $0d915
          55574 => x"00", -- $0d916
          55575 => x"00", -- $0d917
          55576 => x"00", -- $0d918
          55577 => x"00", -- $0d919
          55578 => x"00", -- $0d91a
          55579 => x"00", -- $0d91b
          55580 => x"00", -- $0d91c
          55581 => x"00", -- $0d91d
          55582 => x"00", -- $0d91e
          55583 => x"00", -- $0d91f
          55584 => x"00", -- $0d920
          55585 => x"00", -- $0d921
          55586 => x"00", -- $0d922
          55587 => x"00", -- $0d923
          55588 => x"00", -- $0d924
          55589 => x"00", -- $0d925
          55590 => x"00", -- $0d926
          55591 => x"00", -- $0d927
          55592 => x"00", -- $0d928
          55593 => x"00", -- $0d929
          55594 => x"00", -- $0d92a
          55595 => x"00", -- $0d92b
          55596 => x"00", -- $0d92c
          55597 => x"00", -- $0d92d
          55598 => x"00", -- $0d92e
          55599 => x"00", -- $0d92f
          55600 => x"00", -- $0d930
          55601 => x"00", -- $0d931
          55602 => x"00", -- $0d932
          55603 => x"00", -- $0d933
          55604 => x"00", -- $0d934
          55605 => x"00", -- $0d935
          55606 => x"00", -- $0d936
          55607 => x"00", -- $0d937
          55608 => x"00", -- $0d938
          55609 => x"00", -- $0d939
          55610 => x"00", -- $0d93a
          55611 => x"00", -- $0d93b
          55612 => x"00", -- $0d93c
          55613 => x"00", -- $0d93d
          55614 => x"00", -- $0d93e
          55615 => x"00", -- $0d93f
          55616 => x"00", -- $0d940
          55617 => x"00", -- $0d941
          55618 => x"00", -- $0d942
          55619 => x"00", -- $0d943
          55620 => x"00", -- $0d944
          55621 => x"00", -- $0d945
          55622 => x"00", -- $0d946
          55623 => x"00", -- $0d947
          55624 => x"00", -- $0d948
          55625 => x"00", -- $0d949
          55626 => x"00", -- $0d94a
          55627 => x"00", -- $0d94b
          55628 => x"00", -- $0d94c
          55629 => x"00", -- $0d94d
          55630 => x"00", -- $0d94e
          55631 => x"00", -- $0d94f
          55632 => x"00", -- $0d950
          55633 => x"00", -- $0d951
          55634 => x"00", -- $0d952
          55635 => x"00", -- $0d953
          55636 => x"00", -- $0d954
          55637 => x"00", -- $0d955
          55638 => x"00", -- $0d956
          55639 => x"00", -- $0d957
          55640 => x"00", -- $0d958
          55641 => x"00", -- $0d959
          55642 => x"00", -- $0d95a
          55643 => x"00", -- $0d95b
          55644 => x"00", -- $0d95c
          55645 => x"00", -- $0d95d
          55646 => x"00", -- $0d95e
          55647 => x"00", -- $0d95f
          55648 => x"00", -- $0d960
          55649 => x"00", -- $0d961
          55650 => x"00", -- $0d962
          55651 => x"00", -- $0d963
          55652 => x"00", -- $0d964
          55653 => x"00", -- $0d965
          55654 => x"00", -- $0d966
          55655 => x"00", -- $0d967
          55656 => x"00", -- $0d968
          55657 => x"00", -- $0d969
          55658 => x"00", -- $0d96a
          55659 => x"00", -- $0d96b
          55660 => x"00", -- $0d96c
          55661 => x"00", -- $0d96d
          55662 => x"00", -- $0d96e
          55663 => x"00", -- $0d96f
          55664 => x"00", -- $0d970
          55665 => x"00", -- $0d971
          55666 => x"00", -- $0d972
          55667 => x"00", -- $0d973
          55668 => x"00", -- $0d974
          55669 => x"00", -- $0d975
          55670 => x"00", -- $0d976
          55671 => x"00", -- $0d977
          55672 => x"00", -- $0d978
          55673 => x"00", -- $0d979
          55674 => x"00", -- $0d97a
          55675 => x"00", -- $0d97b
          55676 => x"00", -- $0d97c
          55677 => x"00", -- $0d97d
          55678 => x"00", -- $0d97e
          55679 => x"00", -- $0d97f
          55680 => x"00", -- $0d980
          55681 => x"00", -- $0d981
          55682 => x"00", -- $0d982
          55683 => x"00", -- $0d983
          55684 => x"00", -- $0d984
          55685 => x"00", -- $0d985
          55686 => x"00", -- $0d986
          55687 => x"00", -- $0d987
          55688 => x"00", -- $0d988
          55689 => x"00", -- $0d989
          55690 => x"00", -- $0d98a
          55691 => x"00", -- $0d98b
          55692 => x"00", -- $0d98c
          55693 => x"00", -- $0d98d
          55694 => x"00", -- $0d98e
          55695 => x"00", -- $0d98f
          55696 => x"00", -- $0d990
          55697 => x"00", -- $0d991
          55698 => x"00", -- $0d992
          55699 => x"00", -- $0d993
          55700 => x"00", -- $0d994
          55701 => x"00", -- $0d995
          55702 => x"00", -- $0d996
          55703 => x"00", -- $0d997
          55704 => x"00", -- $0d998
          55705 => x"00", -- $0d999
          55706 => x"00", -- $0d99a
          55707 => x"00", -- $0d99b
          55708 => x"00", -- $0d99c
          55709 => x"00", -- $0d99d
          55710 => x"00", -- $0d99e
          55711 => x"00", -- $0d99f
          55712 => x"00", -- $0d9a0
          55713 => x"00", -- $0d9a1
          55714 => x"00", -- $0d9a2
          55715 => x"00", -- $0d9a3
          55716 => x"00", -- $0d9a4
          55717 => x"00", -- $0d9a5
          55718 => x"00", -- $0d9a6
          55719 => x"00", -- $0d9a7
          55720 => x"00", -- $0d9a8
          55721 => x"00", -- $0d9a9
          55722 => x"00", -- $0d9aa
          55723 => x"00", -- $0d9ab
          55724 => x"00", -- $0d9ac
          55725 => x"00", -- $0d9ad
          55726 => x"00", -- $0d9ae
          55727 => x"00", -- $0d9af
          55728 => x"00", -- $0d9b0
          55729 => x"00", -- $0d9b1
          55730 => x"00", -- $0d9b2
          55731 => x"00", -- $0d9b3
          55732 => x"00", -- $0d9b4
          55733 => x"00", -- $0d9b5
          55734 => x"00", -- $0d9b6
          55735 => x"00", -- $0d9b7
          55736 => x"00", -- $0d9b8
          55737 => x"00", -- $0d9b9
          55738 => x"00", -- $0d9ba
          55739 => x"00", -- $0d9bb
          55740 => x"00", -- $0d9bc
          55741 => x"00", -- $0d9bd
          55742 => x"00", -- $0d9be
          55743 => x"00", -- $0d9bf
          55744 => x"00", -- $0d9c0
          55745 => x"00", -- $0d9c1
          55746 => x"00", -- $0d9c2
          55747 => x"00", -- $0d9c3
          55748 => x"00", -- $0d9c4
          55749 => x"00", -- $0d9c5
          55750 => x"00", -- $0d9c6
          55751 => x"00", -- $0d9c7
          55752 => x"00", -- $0d9c8
          55753 => x"00", -- $0d9c9
          55754 => x"00", -- $0d9ca
          55755 => x"00", -- $0d9cb
          55756 => x"00", -- $0d9cc
          55757 => x"00", -- $0d9cd
          55758 => x"00", -- $0d9ce
          55759 => x"00", -- $0d9cf
          55760 => x"00", -- $0d9d0
          55761 => x"00", -- $0d9d1
          55762 => x"00", -- $0d9d2
          55763 => x"00", -- $0d9d3
          55764 => x"00", -- $0d9d4
          55765 => x"00", -- $0d9d5
          55766 => x"00", -- $0d9d6
          55767 => x"00", -- $0d9d7
          55768 => x"00", -- $0d9d8
          55769 => x"00", -- $0d9d9
          55770 => x"00", -- $0d9da
          55771 => x"00", -- $0d9db
          55772 => x"00", -- $0d9dc
          55773 => x"00", -- $0d9dd
          55774 => x"00", -- $0d9de
          55775 => x"00", -- $0d9df
          55776 => x"00", -- $0d9e0
          55777 => x"00", -- $0d9e1
          55778 => x"00", -- $0d9e2
          55779 => x"00", -- $0d9e3
          55780 => x"00", -- $0d9e4
          55781 => x"00", -- $0d9e5
          55782 => x"00", -- $0d9e6
          55783 => x"00", -- $0d9e7
          55784 => x"00", -- $0d9e8
          55785 => x"00", -- $0d9e9
          55786 => x"00", -- $0d9ea
          55787 => x"00", -- $0d9eb
          55788 => x"00", -- $0d9ec
          55789 => x"00", -- $0d9ed
          55790 => x"00", -- $0d9ee
          55791 => x"00", -- $0d9ef
          55792 => x"00", -- $0d9f0
          55793 => x"00", -- $0d9f1
          55794 => x"00", -- $0d9f2
          55795 => x"00", -- $0d9f3
          55796 => x"00", -- $0d9f4
          55797 => x"00", -- $0d9f5
          55798 => x"00", -- $0d9f6
          55799 => x"00", -- $0d9f7
          55800 => x"00", -- $0d9f8
          55801 => x"00", -- $0d9f9
          55802 => x"00", -- $0d9fa
          55803 => x"00", -- $0d9fb
          55804 => x"00", -- $0d9fc
          55805 => x"00", -- $0d9fd
          55806 => x"00", -- $0d9fe
          55807 => x"00", -- $0d9ff
          55808 => x"00", -- $0da00
          55809 => x"00", -- $0da01
          55810 => x"00", -- $0da02
          55811 => x"00", -- $0da03
          55812 => x"00", -- $0da04
          55813 => x"00", -- $0da05
          55814 => x"00", -- $0da06
          55815 => x"00", -- $0da07
          55816 => x"00", -- $0da08
          55817 => x"00", -- $0da09
          55818 => x"00", -- $0da0a
          55819 => x"00", -- $0da0b
          55820 => x"00", -- $0da0c
          55821 => x"00", -- $0da0d
          55822 => x"00", -- $0da0e
          55823 => x"00", -- $0da0f
          55824 => x"00", -- $0da10
          55825 => x"00", -- $0da11
          55826 => x"00", -- $0da12
          55827 => x"00", -- $0da13
          55828 => x"00", -- $0da14
          55829 => x"00", -- $0da15
          55830 => x"00", -- $0da16
          55831 => x"00", -- $0da17
          55832 => x"00", -- $0da18
          55833 => x"00", -- $0da19
          55834 => x"00", -- $0da1a
          55835 => x"00", -- $0da1b
          55836 => x"00", -- $0da1c
          55837 => x"00", -- $0da1d
          55838 => x"00", -- $0da1e
          55839 => x"00", -- $0da1f
          55840 => x"00", -- $0da20
          55841 => x"00", -- $0da21
          55842 => x"00", -- $0da22
          55843 => x"00", -- $0da23
          55844 => x"00", -- $0da24
          55845 => x"00", -- $0da25
          55846 => x"00", -- $0da26
          55847 => x"00", -- $0da27
          55848 => x"00", -- $0da28
          55849 => x"00", -- $0da29
          55850 => x"00", -- $0da2a
          55851 => x"00", -- $0da2b
          55852 => x"00", -- $0da2c
          55853 => x"00", -- $0da2d
          55854 => x"00", -- $0da2e
          55855 => x"00", -- $0da2f
          55856 => x"00", -- $0da30
          55857 => x"00", -- $0da31
          55858 => x"00", -- $0da32
          55859 => x"00", -- $0da33
          55860 => x"00", -- $0da34
          55861 => x"00", -- $0da35
          55862 => x"00", -- $0da36
          55863 => x"00", -- $0da37
          55864 => x"00", -- $0da38
          55865 => x"00", -- $0da39
          55866 => x"00", -- $0da3a
          55867 => x"00", -- $0da3b
          55868 => x"00", -- $0da3c
          55869 => x"00", -- $0da3d
          55870 => x"00", -- $0da3e
          55871 => x"00", -- $0da3f
          55872 => x"00", -- $0da40
          55873 => x"00", -- $0da41
          55874 => x"00", -- $0da42
          55875 => x"00", -- $0da43
          55876 => x"00", -- $0da44
          55877 => x"00", -- $0da45
          55878 => x"00", -- $0da46
          55879 => x"00", -- $0da47
          55880 => x"00", -- $0da48
          55881 => x"00", -- $0da49
          55882 => x"00", -- $0da4a
          55883 => x"00", -- $0da4b
          55884 => x"00", -- $0da4c
          55885 => x"00", -- $0da4d
          55886 => x"00", -- $0da4e
          55887 => x"00", -- $0da4f
          55888 => x"00", -- $0da50
          55889 => x"00", -- $0da51
          55890 => x"00", -- $0da52
          55891 => x"00", -- $0da53
          55892 => x"00", -- $0da54
          55893 => x"00", -- $0da55
          55894 => x"00", -- $0da56
          55895 => x"00", -- $0da57
          55896 => x"00", -- $0da58
          55897 => x"00", -- $0da59
          55898 => x"00", -- $0da5a
          55899 => x"00", -- $0da5b
          55900 => x"00", -- $0da5c
          55901 => x"00", -- $0da5d
          55902 => x"00", -- $0da5e
          55903 => x"00", -- $0da5f
          55904 => x"00", -- $0da60
          55905 => x"00", -- $0da61
          55906 => x"00", -- $0da62
          55907 => x"00", -- $0da63
          55908 => x"00", -- $0da64
          55909 => x"00", -- $0da65
          55910 => x"00", -- $0da66
          55911 => x"00", -- $0da67
          55912 => x"00", -- $0da68
          55913 => x"00", -- $0da69
          55914 => x"00", -- $0da6a
          55915 => x"00", -- $0da6b
          55916 => x"00", -- $0da6c
          55917 => x"00", -- $0da6d
          55918 => x"00", -- $0da6e
          55919 => x"00", -- $0da6f
          55920 => x"00", -- $0da70
          55921 => x"00", -- $0da71
          55922 => x"00", -- $0da72
          55923 => x"00", -- $0da73
          55924 => x"00", -- $0da74
          55925 => x"00", -- $0da75
          55926 => x"00", -- $0da76
          55927 => x"00", -- $0da77
          55928 => x"00", -- $0da78
          55929 => x"00", -- $0da79
          55930 => x"00", -- $0da7a
          55931 => x"00", -- $0da7b
          55932 => x"00", -- $0da7c
          55933 => x"00", -- $0da7d
          55934 => x"00", -- $0da7e
          55935 => x"00", -- $0da7f
          55936 => x"00", -- $0da80
          55937 => x"00", -- $0da81
          55938 => x"00", -- $0da82
          55939 => x"00", -- $0da83
          55940 => x"00", -- $0da84
          55941 => x"00", -- $0da85
          55942 => x"00", -- $0da86
          55943 => x"00", -- $0da87
          55944 => x"00", -- $0da88
          55945 => x"00", -- $0da89
          55946 => x"00", -- $0da8a
          55947 => x"00", -- $0da8b
          55948 => x"00", -- $0da8c
          55949 => x"00", -- $0da8d
          55950 => x"00", -- $0da8e
          55951 => x"00", -- $0da8f
          55952 => x"00", -- $0da90
          55953 => x"00", -- $0da91
          55954 => x"00", -- $0da92
          55955 => x"00", -- $0da93
          55956 => x"00", -- $0da94
          55957 => x"00", -- $0da95
          55958 => x"00", -- $0da96
          55959 => x"00", -- $0da97
          55960 => x"00", -- $0da98
          55961 => x"00", -- $0da99
          55962 => x"00", -- $0da9a
          55963 => x"00", -- $0da9b
          55964 => x"00", -- $0da9c
          55965 => x"00", -- $0da9d
          55966 => x"00", -- $0da9e
          55967 => x"00", -- $0da9f
          55968 => x"00", -- $0daa0
          55969 => x"00", -- $0daa1
          55970 => x"00", -- $0daa2
          55971 => x"00", -- $0daa3
          55972 => x"00", -- $0daa4
          55973 => x"00", -- $0daa5
          55974 => x"00", -- $0daa6
          55975 => x"00", -- $0daa7
          55976 => x"00", -- $0daa8
          55977 => x"00", -- $0daa9
          55978 => x"00", -- $0daaa
          55979 => x"00", -- $0daab
          55980 => x"00", -- $0daac
          55981 => x"00", -- $0daad
          55982 => x"00", -- $0daae
          55983 => x"00", -- $0daaf
          55984 => x"00", -- $0dab0
          55985 => x"00", -- $0dab1
          55986 => x"00", -- $0dab2
          55987 => x"00", -- $0dab3
          55988 => x"00", -- $0dab4
          55989 => x"00", -- $0dab5
          55990 => x"00", -- $0dab6
          55991 => x"00", -- $0dab7
          55992 => x"00", -- $0dab8
          55993 => x"00", -- $0dab9
          55994 => x"00", -- $0daba
          55995 => x"00", -- $0dabb
          55996 => x"00", -- $0dabc
          55997 => x"00", -- $0dabd
          55998 => x"00", -- $0dabe
          55999 => x"00", -- $0dabf
          56000 => x"00", -- $0dac0
          56001 => x"00", -- $0dac1
          56002 => x"00", -- $0dac2
          56003 => x"00", -- $0dac3
          56004 => x"00", -- $0dac4
          56005 => x"00", -- $0dac5
          56006 => x"00", -- $0dac6
          56007 => x"00", -- $0dac7
          56008 => x"00", -- $0dac8
          56009 => x"00", -- $0dac9
          56010 => x"00", -- $0daca
          56011 => x"00", -- $0dacb
          56012 => x"00", -- $0dacc
          56013 => x"00", -- $0dacd
          56014 => x"00", -- $0dace
          56015 => x"00", -- $0dacf
          56016 => x"00", -- $0dad0
          56017 => x"00", -- $0dad1
          56018 => x"00", -- $0dad2
          56019 => x"00", -- $0dad3
          56020 => x"00", -- $0dad4
          56021 => x"00", -- $0dad5
          56022 => x"00", -- $0dad6
          56023 => x"00", -- $0dad7
          56024 => x"00", -- $0dad8
          56025 => x"00", -- $0dad9
          56026 => x"00", -- $0dada
          56027 => x"00", -- $0dadb
          56028 => x"00", -- $0dadc
          56029 => x"00", -- $0dadd
          56030 => x"00", -- $0dade
          56031 => x"00", -- $0dadf
          56032 => x"00", -- $0dae0
          56033 => x"00", -- $0dae1
          56034 => x"00", -- $0dae2
          56035 => x"00", -- $0dae3
          56036 => x"00", -- $0dae4
          56037 => x"00", -- $0dae5
          56038 => x"00", -- $0dae6
          56039 => x"00", -- $0dae7
          56040 => x"00", -- $0dae8
          56041 => x"00", -- $0dae9
          56042 => x"00", -- $0daea
          56043 => x"00", -- $0daeb
          56044 => x"00", -- $0daec
          56045 => x"00", -- $0daed
          56046 => x"00", -- $0daee
          56047 => x"00", -- $0daef
          56048 => x"00", -- $0daf0
          56049 => x"00", -- $0daf1
          56050 => x"00", -- $0daf2
          56051 => x"00", -- $0daf3
          56052 => x"00", -- $0daf4
          56053 => x"00", -- $0daf5
          56054 => x"00", -- $0daf6
          56055 => x"00", -- $0daf7
          56056 => x"00", -- $0daf8
          56057 => x"00", -- $0daf9
          56058 => x"00", -- $0dafa
          56059 => x"00", -- $0dafb
          56060 => x"00", -- $0dafc
          56061 => x"00", -- $0dafd
          56062 => x"00", -- $0dafe
          56063 => x"00", -- $0daff
          56064 => x"00", -- $0db00
          56065 => x"00", -- $0db01
          56066 => x"00", -- $0db02
          56067 => x"00", -- $0db03
          56068 => x"00", -- $0db04
          56069 => x"00", -- $0db05
          56070 => x"00", -- $0db06
          56071 => x"00", -- $0db07
          56072 => x"00", -- $0db08
          56073 => x"00", -- $0db09
          56074 => x"00", -- $0db0a
          56075 => x"00", -- $0db0b
          56076 => x"00", -- $0db0c
          56077 => x"00", -- $0db0d
          56078 => x"00", -- $0db0e
          56079 => x"00", -- $0db0f
          56080 => x"00", -- $0db10
          56081 => x"00", -- $0db11
          56082 => x"00", -- $0db12
          56083 => x"00", -- $0db13
          56084 => x"00", -- $0db14
          56085 => x"00", -- $0db15
          56086 => x"00", -- $0db16
          56087 => x"00", -- $0db17
          56088 => x"00", -- $0db18
          56089 => x"00", -- $0db19
          56090 => x"00", -- $0db1a
          56091 => x"00", -- $0db1b
          56092 => x"00", -- $0db1c
          56093 => x"00", -- $0db1d
          56094 => x"00", -- $0db1e
          56095 => x"00", -- $0db1f
          56096 => x"00", -- $0db20
          56097 => x"00", -- $0db21
          56098 => x"00", -- $0db22
          56099 => x"00", -- $0db23
          56100 => x"00", -- $0db24
          56101 => x"00", -- $0db25
          56102 => x"00", -- $0db26
          56103 => x"00", -- $0db27
          56104 => x"00", -- $0db28
          56105 => x"00", -- $0db29
          56106 => x"00", -- $0db2a
          56107 => x"00", -- $0db2b
          56108 => x"00", -- $0db2c
          56109 => x"00", -- $0db2d
          56110 => x"00", -- $0db2e
          56111 => x"00", -- $0db2f
          56112 => x"00", -- $0db30
          56113 => x"00", -- $0db31
          56114 => x"00", -- $0db32
          56115 => x"00", -- $0db33
          56116 => x"00", -- $0db34
          56117 => x"00", -- $0db35
          56118 => x"00", -- $0db36
          56119 => x"00", -- $0db37
          56120 => x"00", -- $0db38
          56121 => x"00", -- $0db39
          56122 => x"00", -- $0db3a
          56123 => x"00", -- $0db3b
          56124 => x"00", -- $0db3c
          56125 => x"00", -- $0db3d
          56126 => x"00", -- $0db3e
          56127 => x"00", -- $0db3f
          56128 => x"00", -- $0db40
          56129 => x"00", -- $0db41
          56130 => x"00", -- $0db42
          56131 => x"00", -- $0db43
          56132 => x"00", -- $0db44
          56133 => x"00", -- $0db45
          56134 => x"00", -- $0db46
          56135 => x"00", -- $0db47
          56136 => x"00", -- $0db48
          56137 => x"00", -- $0db49
          56138 => x"00", -- $0db4a
          56139 => x"00", -- $0db4b
          56140 => x"00", -- $0db4c
          56141 => x"00", -- $0db4d
          56142 => x"00", -- $0db4e
          56143 => x"00", -- $0db4f
          56144 => x"00", -- $0db50
          56145 => x"00", -- $0db51
          56146 => x"00", -- $0db52
          56147 => x"00", -- $0db53
          56148 => x"00", -- $0db54
          56149 => x"00", -- $0db55
          56150 => x"00", -- $0db56
          56151 => x"00", -- $0db57
          56152 => x"00", -- $0db58
          56153 => x"00", -- $0db59
          56154 => x"00", -- $0db5a
          56155 => x"00", -- $0db5b
          56156 => x"00", -- $0db5c
          56157 => x"00", -- $0db5d
          56158 => x"00", -- $0db5e
          56159 => x"00", -- $0db5f
          56160 => x"00", -- $0db60
          56161 => x"00", -- $0db61
          56162 => x"00", -- $0db62
          56163 => x"00", -- $0db63
          56164 => x"00", -- $0db64
          56165 => x"00", -- $0db65
          56166 => x"00", -- $0db66
          56167 => x"00", -- $0db67
          56168 => x"00", -- $0db68
          56169 => x"00", -- $0db69
          56170 => x"00", -- $0db6a
          56171 => x"00", -- $0db6b
          56172 => x"00", -- $0db6c
          56173 => x"00", -- $0db6d
          56174 => x"00", -- $0db6e
          56175 => x"00", -- $0db6f
          56176 => x"00", -- $0db70
          56177 => x"00", -- $0db71
          56178 => x"00", -- $0db72
          56179 => x"00", -- $0db73
          56180 => x"00", -- $0db74
          56181 => x"00", -- $0db75
          56182 => x"00", -- $0db76
          56183 => x"00", -- $0db77
          56184 => x"00", -- $0db78
          56185 => x"00", -- $0db79
          56186 => x"00", -- $0db7a
          56187 => x"00", -- $0db7b
          56188 => x"00", -- $0db7c
          56189 => x"00", -- $0db7d
          56190 => x"00", -- $0db7e
          56191 => x"00", -- $0db7f
          56192 => x"00", -- $0db80
          56193 => x"00", -- $0db81
          56194 => x"00", -- $0db82
          56195 => x"00", -- $0db83
          56196 => x"00", -- $0db84
          56197 => x"00", -- $0db85
          56198 => x"00", -- $0db86
          56199 => x"00", -- $0db87
          56200 => x"00", -- $0db88
          56201 => x"00", -- $0db89
          56202 => x"00", -- $0db8a
          56203 => x"00", -- $0db8b
          56204 => x"00", -- $0db8c
          56205 => x"00", -- $0db8d
          56206 => x"00", -- $0db8e
          56207 => x"00", -- $0db8f
          56208 => x"00", -- $0db90
          56209 => x"00", -- $0db91
          56210 => x"00", -- $0db92
          56211 => x"00", -- $0db93
          56212 => x"00", -- $0db94
          56213 => x"00", -- $0db95
          56214 => x"00", -- $0db96
          56215 => x"00", -- $0db97
          56216 => x"00", -- $0db98
          56217 => x"00", -- $0db99
          56218 => x"00", -- $0db9a
          56219 => x"00", -- $0db9b
          56220 => x"00", -- $0db9c
          56221 => x"00", -- $0db9d
          56222 => x"00", -- $0db9e
          56223 => x"00", -- $0db9f
          56224 => x"00", -- $0dba0
          56225 => x"00", -- $0dba1
          56226 => x"00", -- $0dba2
          56227 => x"00", -- $0dba3
          56228 => x"00", -- $0dba4
          56229 => x"00", -- $0dba5
          56230 => x"00", -- $0dba6
          56231 => x"00", -- $0dba7
          56232 => x"00", -- $0dba8
          56233 => x"00", -- $0dba9
          56234 => x"00", -- $0dbaa
          56235 => x"00", -- $0dbab
          56236 => x"00", -- $0dbac
          56237 => x"00", -- $0dbad
          56238 => x"00", -- $0dbae
          56239 => x"00", -- $0dbaf
          56240 => x"00", -- $0dbb0
          56241 => x"00", -- $0dbb1
          56242 => x"00", -- $0dbb2
          56243 => x"00", -- $0dbb3
          56244 => x"00", -- $0dbb4
          56245 => x"00", -- $0dbb5
          56246 => x"00", -- $0dbb6
          56247 => x"00", -- $0dbb7
          56248 => x"00", -- $0dbb8
          56249 => x"00", -- $0dbb9
          56250 => x"00", -- $0dbba
          56251 => x"00", -- $0dbbb
          56252 => x"00", -- $0dbbc
          56253 => x"00", -- $0dbbd
          56254 => x"00", -- $0dbbe
          56255 => x"00", -- $0dbbf
          56256 => x"00", -- $0dbc0
          56257 => x"00", -- $0dbc1
          56258 => x"00", -- $0dbc2
          56259 => x"00", -- $0dbc3
          56260 => x"00", -- $0dbc4
          56261 => x"00", -- $0dbc5
          56262 => x"00", -- $0dbc6
          56263 => x"00", -- $0dbc7
          56264 => x"00", -- $0dbc8
          56265 => x"00", -- $0dbc9
          56266 => x"00", -- $0dbca
          56267 => x"00", -- $0dbcb
          56268 => x"00", -- $0dbcc
          56269 => x"00", -- $0dbcd
          56270 => x"00", -- $0dbce
          56271 => x"00", -- $0dbcf
          56272 => x"00", -- $0dbd0
          56273 => x"00", -- $0dbd1
          56274 => x"00", -- $0dbd2
          56275 => x"00", -- $0dbd3
          56276 => x"00", -- $0dbd4
          56277 => x"00", -- $0dbd5
          56278 => x"00", -- $0dbd6
          56279 => x"00", -- $0dbd7
          56280 => x"00", -- $0dbd8
          56281 => x"00", -- $0dbd9
          56282 => x"00", -- $0dbda
          56283 => x"00", -- $0dbdb
          56284 => x"00", -- $0dbdc
          56285 => x"00", -- $0dbdd
          56286 => x"00", -- $0dbde
          56287 => x"00", -- $0dbdf
          56288 => x"00", -- $0dbe0
          56289 => x"00", -- $0dbe1
          56290 => x"00", -- $0dbe2
          56291 => x"00", -- $0dbe3
          56292 => x"00", -- $0dbe4
          56293 => x"00", -- $0dbe5
          56294 => x"00", -- $0dbe6
          56295 => x"00", -- $0dbe7
          56296 => x"00", -- $0dbe8
          56297 => x"00", -- $0dbe9
          56298 => x"00", -- $0dbea
          56299 => x"00", -- $0dbeb
          56300 => x"00", -- $0dbec
          56301 => x"00", -- $0dbed
          56302 => x"00", -- $0dbee
          56303 => x"00", -- $0dbef
          56304 => x"00", -- $0dbf0
          56305 => x"00", -- $0dbf1
          56306 => x"00", -- $0dbf2
          56307 => x"00", -- $0dbf3
          56308 => x"00", -- $0dbf4
          56309 => x"00", -- $0dbf5
          56310 => x"00", -- $0dbf6
          56311 => x"00", -- $0dbf7
          56312 => x"00", -- $0dbf8
          56313 => x"00", -- $0dbf9
          56314 => x"00", -- $0dbfa
          56315 => x"00", -- $0dbfb
          56316 => x"00", -- $0dbfc
          56317 => x"00", -- $0dbfd
          56318 => x"00", -- $0dbfe
          56319 => x"00", -- $0dbff
          56320 => x"00", -- $0dc00
          56321 => x"00", -- $0dc01
          56322 => x"00", -- $0dc02
          56323 => x"00", -- $0dc03
          56324 => x"00", -- $0dc04
          56325 => x"00", -- $0dc05
          56326 => x"00", -- $0dc06
          56327 => x"00", -- $0dc07
          56328 => x"00", -- $0dc08
          56329 => x"00", -- $0dc09
          56330 => x"00", -- $0dc0a
          56331 => x"00", -- $0dc0b
          56332 => x"00", -- $0dc0c
          56333 => x"00", -- $0dc0d
          56334 => x"00", -- $0dc0e
          56335 => x"00", -- $0dc0f
          56336 => x"00", -- $0dc10
          56337 => x"00", -- $0dc11
          56338 => x"00", -- $0dc12
          56339 => x"00", -- $0dc13
          56340 => x"00", -- $0dc14
          56341 => x"00", -- $0dc15
          56342 => x"00", -- $0dc16
          56343 => x"00", -- $0dc17
          56344 => x"00", -- $0dc18
          56345 => x"00", -- $0dc19
          56346 => x"00", -- $0dc1a
          56347 => x"00", -- $0dc1b
          56348 => x"00", -- $0dc1c
          56349 => x"00", -- $0dc1d
          56350 => x"00", -- $0dc1e
          56351 => x"00", -- $0dc1f
          56352 => x"00", -- $0dc20
          56353 => x"00", -- $0dc21
          56354 => x"00", -- $0dc22
          56355 => x"00", -- $0dc23
          56356 => x"00", -- $0dc24
          56357 => x"00", -- $0dc25
          56358 => x"00", -- $0dc26
          56359 => x"00", -- $0dc27
          56360 => x"00", -- $0dc28
          56361 => x"00", -- $0dc29
          56362 => x"00", -- $0dc2a
          56363 => x"00", -- $0dc2b
          56364 => x"00", -- $0dc2c
          56365 => x"00", -- $0dc2d
          56366 => x"00", -- $0dc2e
          56367 => x"00", -- $0dc2f
          56368 => x"00", -- $0dc30
          56369 => x"00", -- $0dc31
          56370 => x"00", -- $0dc32
          56371 => x"00", -- $0dc33
          56372 => x"00", -- $0dc34
          56373 => x"00", -- $0dc35
          56374 => x"00", -- $0dc36
          56375 => x"00", -- $0dc37
          56376 => x"00", -- $0dc38
          56377 => x"00", -- $0dc39
          56378 => x"00", -- $0dc3a
          56379 => x"00", -- $0dc3b
          56380 => x"00", -- $0dc3c
          56381 => x"00", -- $0dc3d
          56382 => x"00", -- $0dc3e
          56383 => x"00", -- $0dc3f
          56384 => x"00", -- $0dc40
          56385 => x"00", -- $0dc41
          56386 => x"00", -- $0dc42
          56387 => x"00", -- $0dc43
          56388 => x"00", -- $0dc44
          56389 => x"00", -- $0dc45
          56390 => x"00", -- $0dc46
          56391 => x"00", -- $0dc47
          56392 => x"00", -- $0dc48
          56393 => x"00", -- $0dc49
          56394 => x"00", -- $0dc4a
          56395 => x"00", -- $0dc4b
          56396 => x"00", -- $0dc4c
          56397 => x"00", -- $0dc4d
          56398 => x"00", -- $0dc4e
          56399 => x"00", -- $0dc4f
          56400 => x"00", -- $0dc50
          56401 => x"00", -- $0dc51
          56402 => x"00", -- $0dc52
          56403 => x"00", -- $0dc53
          56404 => x"00", -- $0dc54
          56405 => x"00", -- $0dc55
          56406 => x"00", -- $0dc56
          56407 => x"00", -- $0dc57
          56408 => x"00", -- $0dc58
          56409 => x"00", -- $0dc59
          56410 => x"00", -- $0dc5a
          56411 => x"00", -- $0dc5b
          56412 => x"00", -- $0dc5c
          56413 => x"00", -- $0dc5d
          56414 => x"00", -- $0dc5e
          56415 => x"00", -- $0dc5f
          56416 => x"00", -- $0dc60
          56417 => x"00", -- $0dc61
          56418 => x"00", -- $0dc62
          56419 => x"00", -- $0dc63
          56420 => x"00", -- $0dc64
          56421 => x"00", -- $0dc65
          56422 => x"00", -- $0dc66
          56423 => x"00", -- $0dc67
          56424 => x"00", -- $0dc68
          56425 => x"00", -- $0dc69
          56426 => x"00", -- $0dc6a
          56427 => x"00", -- $0dc6b
          56428 => x"00", -- $0dc6c
          56429 => x"00", -- $0dc6d
          56430 => x"00", -- $0dc6e
          56431 => x"00", -- $0dc6f
          56432 => x"00", -- $0dc70
          56433 => x"00", -- $0dc71
          56434 => x"00", -- $0dc72
          56435 => x"00", -- $0dc73
          56436 => x"00", -- $0dc74
          56437 => x"00", -- $0dc75
          56438 => x"00", -- $0dc76
          56439 => x"00", -- $0dc77
          56440 => x"00", -- $0dc78
          56441 => x"00", -- $0dc79
          56442 => x"00", -- $0dc7a
          56443 => x"00", -- $0dc7b
          56444 => x"00", -- $0dc7c
          56445 => x"00", -- $0dc7d
          56446 => x"00", -- $0dc7e
          56447 => x"00", -- $0dc7f
          56448 => x"00", -- $0dc80
          56449 => x"00", -- $0dc81
          56450 => x"00", -- $0dc82
          56451 => x"00", -- $0dc83
          56452 => x"00", -- $0dc84
          56453 => x"00", -- $0dc85
          56454 => x"00", -- $0dc86
          56455 => x"00", -- $0dc87
          56456 => x"00", -- $0dc88
          56457 => x"00", -- $0dc89
          56458 => x"00", -- $0dc8a
          56459 => x"00", -- $0dc8b
          56460 => x"00", -- $0dc8c
          56461 => x"00", -- $0dc8d
          56462 => x"00", -- $0dc8e
          56463 => x"00", -- $0dc8f
          56464 => x"00", -- $0dc90
          56465 => x"00", -- $0dc91
          56466 => x"00", -- $0dc92
          56467 => x"00", -- $0dc93
          56468 => x"00", -- $0dc94
          56469 => x"00", -- $0dc95
          56470 => x"00", -- $0dc96
          56471 => x"00", -- $0dc97
          56472 => x"00", -- $0dc98
          56473 => x"00", -- $0dc99
          56474 => x"00", -- $0dc9a
          56475 => x"00", -- $0dc9b
          56476 => x"00", -- $0dc9c
          56477 => x"00", -- $0dc9d
          56478 => x"00", -- $0dc9e
          56479 => x"00", -- $0dc9f
          56480 => x"00", -- $0dca0
          56481 => x"00", -- $0dca1
          56482 => x"00", -- $0dca2
          56483 => x"00", -- $0dca3
          56484 => x"00", -- $0dca4
          56485 => x"00", -- $0dca5
          56486 => x"00", -- $0dca6
          56487 => x"00", -- $0dca7
          56488 => x"00", -- $0dca8
          56489 => x"00", -- $0dca9
          56490 => x"00", -- $0dcaa
          56491 => x"00", -- $0dcab
          56492 => x"00", -- $0dcac
          56493 => x"00", -- $0dcad
          56494 => x"00", -- $0dcae
          56495 => x"00", -- $0dcaf
          56496 => x"00", -- $0dcb0
          56497 => x"00", -- $0dcb1
          56498 => x"00", -- $0dcb2
          56499 => x"00", -- $0dcb3
          56500 => x"00", -- $0dcb4
          56501 => x"00", -- $0dcb5
          56502 => x"00", -- $0dcb6
          56503 => x"00", -- $0dcb7
          56504 => x"00", -- $0dcb8
          56505 => x"00", -- $0dcb9
          56506 => x"00", -- $0dcba
          56507 => x"00", -- $0dcbb
          56508 => x"00", -- $0dcbc
          56509 => x"00", -- $0dcbd
          56510 => x"00", -- $0dcbe
          56511 => x"00", -- $0dcbf
          56512 => x"00", -- $0dcc0
          56513 => x"00", -- $0dcc1
          56514 => x"00", -- $0dcc2
          56515 => x"00", -- $0dcc3
          56516 => x"00", -- $0dcc4
          56517 => x"00", -- $0dcc5
          56518 => x"00", -- $0dcc6
          56519 => x"00", -- $0dcc7
          56520 => x"00", -- $0dcc8
          56521 => x"00", -- $0dcc9
          56522 => x"00", -- $0dcca
          56523 => x"00", -- $0dccb
          56524 => x"00", -- $0dccc
          56525 => x"00", -- $0dccd
          56526 => x"00", -- $0dcce
          56527 => x"00", -- $0dccf
          56528 => x"00", -- $0dcd0
          56529 => x"00", -- $0dcd1
          56530 => x"00", -- $0dcd2
          56531 => x"00", -- $0dcd3
          56532 => x"00", -- $0dcd4
          56533 => x"00", -- $0dcd5
          56534 => x"00", -- $0dcd6
          56535 => x"00", -- $0dcd7
          56536 => x"00", -- $0dcd8
          56537 => x"00", -- $0dcd9
          56538 => x"00", -- $0dcda
          56539 => x"00", -- $0dcdb
          56540 => x"00", -- $0dcdc
          56541 => x"00", -- $0dcdd
          56542 => x"00", -- $0dcde
          56543 => x"00", -- $0dcdf
          56544 => x"00", -- $0dce0
          56545 => x"00", -- $0dce1
          56546 => x"00", -- $0dce2
          56547 => x"00", -- $0dce3
          56548 => x"00", -- $0dce4
          56549 => x"00", -- $0dce5
          56550 => x"00", -- $0dce6
          56551 => x"00", -- $0dce7
          56552 => x"00", -- $0dce8
          56553 => x"00", -- $0dce9
          56554 => x"00", -- $0dcea
          56555 => x"00", -- $0dceb
          56556 => x"00", -- $0dcec
          56557 => x"00", -- $0dced
          56558 => x"00", -- $0dcee
          56559 => x"00", -- $0dcef
          56560 => x"00", -- $0dcf0
          56561 => x"00", -- $0dcf1
          56562 => x"00", -- $0dcf2
          56563 => x"00", -- $0dcf3
          56564 => x"00", -- $0dcf4
          56565 => x"00", -- $0dcf5
          56566 => x"00", -- $0dcf6
          56567 => x"00", -- $0dcf7
          56568 => x"00", -- $0dcf8
          56569 => x"00", -- $0dcf9
          56570 => x"00", -- $0dcfa
          56571 => x"00", -- $0dcfb
          56572 => x"00", -- $0dcfc
          56573 => x"00", -- $0dcfd
          56574 => x"00", -- $0dcfe
          56575 => x"00", -- $0dcff
          56576 => x"00", -- $0dd00
          56577 => x"00", -- $0dd01
          56578 => x"00", -- $0dd02
          56579 => x"00", -- $0dd03
          56580 => x"00", -- $0dd04
          56581 => x"00", -- $0dd05
          56582 => x"00", -- $0dd06
          56583 => x"00", -- $0dd07
          56584 => x"00", -- $0dd08
          56585 => x"00", -- $0dd09
          56586 => x"00", -- $0dd0a
          56587 => x"00", -- $0dd0b
          56588 => x"00", -- $0dd0c
          56589 => x"00", -- $0dd0d
          56590 => x"00", -- $0dd0e
          56591 => x"00", -- $0dd0f
          56592 => x"00", -- $0dd10
          56593 => x"00", -- $0dd11
          56594 => x"00", -- $0dd12
          56595 => x"00", -- $0dd13
          56596 => x"00", -- $0dd14
          56597 => x"00", -- $0dd15
          56598 => x"00", -- $0dd16
          56599 => x"00", -- $0dd17
          56600 => x"00", -- $0dd18
          56601 => x"00", -- $0dd19
          56602 => x"00", -- $0dd1a
          56603 => x"00", -- $0dd1b
          56604 => x"00", -- $0dd1c
          56605 => x"00", -- $0dd1d
          56606 => x"00", -- $0dd1e
          56607 => x"00", -- $0dd1f
          56608 => x"00", -- $0dd20
          56609 => x"00", -- $0dd21
          56610 => x"00", -- $0dd22
          56611 => x"00", -- $0dd23
          56612 => x"00", -- $0dd24
          56613 => x"00", -- $0dd25
          56614 => x"00", -- $0dd26
          56615 => x"00", -- $0dd27
          56616 => x"00", -- $0dd28
          56617 => x"00", -- $0dd29
          56618 => x"00", -- $0dd2a
          56619 => x"00", -- $0dd2b
          56620 => x"00", -- $0dd2c
          56621 => x"00", -- $0dd2d
          56622 => x"00", -- $0dd2e
          56623 => x"00", -- $0dd2f
          56624 => x"00", -- $0dd30
          56625 => x"00", -- $0dd31
          56626 => x"00", -- $0dd32
          56627 => x"00", -- $0dd33
          56628 => x"00", -- $0dd34
          56629 => x"00", -- $0dd35
          56630 => x"00", -- $0dd36
          56631 => x"00", -- $0dd37
          56632 => x"00", -- $0dd38
          56633 => x"00", -- $0dd39
          56634 => x"00", -- $0dd3a
          56635 => x"00", -- $0dd3b
          56636 => x"00", -- $0dd3c
          56637 => x"00", -- $0dd3d
          56638 => x"00", -- $0dd3e
          56639 => x"00", -- $0dd3f
          56640 => x"00", -- $0dd40
          56641 => x"00", -- $0dd41
          56642 => x"00", -- $0dd42
          56643 => x"00", -- $0dd43
          56644 => x"00", -- $0dd44
          56645 => x"00", -- $0dd45
          56646 => x"00", -- $0dd46
          56647 => x"00", -- $0dd47
          56648 => x"00", -- $0dd48
          56649 => x"00", -- $0dd49
          56650 => x"00", -- $0dd4a
          56651 => x"00", -- $0dd4b
          56652 => x"00", -- $0dd4c
          56653 => x"00", -- $0dd4d
          56654 => x"00", -- $0dd4e
          56655 => x"00", -- $0dd4f
          56656 => x"00", -- $0dd50
          56657 => x"00", -- $0dd51
          56658 => x"00", -- $0dd52
          56659 => x"00", -- $0dd53
          56660 => x"00", -- $0dd54
          56661 => x"00", -- $0dd55
          56662 => x"00", -- $0dd56
          56663 => x"00", -- $0dd57
          56664 => x"00", -- $0dd58
          56665 => x"00", -- $0dd59
          56666 => x"00", -- $0dd5a
          56667 => x"00", -- $0dd5b
          56668 => x"00", -- $0dd5c
          56669 => x"00", -- $0dd5d
          56670 => x"00", -- $0dd5e
          56671 => x"00", -- $0dd5f
          56672 => x"00", -- $0dd60
          56673 => x"00", -- $0dd61
          56674 => x"00", -- $0dd62
          56675 => x"00", -- $0dd63
          56676 => x"00", -- $0dd64
          56677 => x"00", -- $0dd65
          56678 => x"00", -- $0dd66
          56679 => x"00", -- $0dd67
          56680 => x"00", -- $0dd68
          56681 => x"00", -- $0dd69
          56682 => x"00", -- $0dd6a
          56683 => x"00", -- $0dd6b
          56684 => x"00", -- $0dd6c
          56685 => x"00", -- $0dd6d
          56686 => x"00", -- $0dd6e
          56687 => x"00", -- $0dd6f
          56688 => x"00", -- $0dd70
          56689 => x"00", -- $0dd71
          56690 => x"00", -- $0dd72
          56691 => x"00", -- $0dd73
          56692 => x"00", -- $0dd74
          56693 => x"00", -- $0dd75
          56694 => x"00", -- $0dd76
          56695 => x"00", -- $0dd77
          56696 => x"00", -- $0dd78
          56697 => x"00", -- $0dd79
          56698 => x"00", -- $0dd7a
          56699 => x"00", -- $0dd7b
          56700 => x"00", -- $0dd7c
          56701 => x"00", -- $0dd7d
          56702 => x"00", -- $0dd7e
          56703 => x"00", -- $0dd7f
          56704 => x"00", -- $0dd80
          56705 => x"00", -- $0dd81
          56706 => x"00", -- $0dd82
          56707 => x"00", -- $0dd83
          56708 => x"00", -- $0dd84
          56709 => x"00", -- $0dd85
          56710 => x"00", -- $0dd86
          56711 => x"00", -- $0dd87
          56712 => x"00", -- $0dd88
          56713 => x"00", -- $0dd89
          56714 => x"00", -- $0dd8a
          56715 => x"00", -- $0dd8b
          56716 => x"00", -- $0dd8c
          56717 => x"00", -- $0dd8d
          56718 => x"00", -- $0dd8e
          56719 => x"00", -- $0dd8f
          56720 => x"00", -- $0dd90
          56721 => x"00", -- $0dd91
          56722 => x"00", -- $0dd92
          56723 => x"00", -- $0dd93
          56724 => x"00", -- $0dd94
          56725 => x"00", -- $0dd95
          56726 => x"00", -- $0dd96
          56727 => x"00", -- $0dd97
          56728 => x"00", -- $0dd98
          56729 => x"00", -- $0dd99
          56730 => x"00", -- $0dd9a
          56731 => x"00", -- $0dd9b
          56732 => x"00", -- $0dd9c
          56733 => x"00", -- $0dd9d
          56734 => x"00", -- $0dd9e
          56735 => x"00", -- $0dd9f
          56736 => x"00", -- $0dda0
          56737 => x"00", -- $0dda1
          56738 => x"00", -- $0dda2
          56739 => x"00", -- $0dda3
          56740 => x"00", -- $0dda4
          56741 => x"00", -- $0dda5
          56742 => x"00", -- $0dda6
          56743 => x"00", -- $0dda7
          56744 => x"00", -- $0dda8
          56745 => x"00", -- $0dda9
          56746 => x"00", -- $0ddaa
          56747 => x"00", -- $0ddab
          56748 => x"00", -- $0ddac
          56749 => x"00", -- $0ddad
          56750 => x"00", -- $0ddae
          56751 => x"00", -- $0ddaf
          56752 => x"00", -- $0ddb0
          56753 => x"00", -- $0ddb1
          56754 => x"00", -- $0ddb2
          56755 => x"00", -- $0ddb3
          56756 => x"00", -- $0ddb4
          56757 => x"00", -- $0ddb5
          56758 => x"00", -- $0ddb6
          56759 => x"00", -- $0ddb7
          56760 => x"00", -- $0ddb8
          56761 => x"00", -- $0ddb9
          56762 => x"00", -- $0ddba
          56763 => x"00", -- $0ddbb
          56764 => x"00", -- $0ddbc
          56765 => x"00", -- $0ddbd
          56766 => x"00", -- $0ddbe
          56767 => x"00", -- $0ddbf
          56768 => x"00", -- $0ddc0
          56769 => x"00", -- $0ddc1
          56770 => x"00", -- $0ddc2
          56771 => x"00", -- $0ddc3
          56772 => x"00", -- $0ddc4
          56773 => x"00", -- $0ddc5
          56774 => x"00", -- $0ddc6
          56775 => x"00", -- $0ddc7
          56776 => x"00", -- $0ddc8
          56777 => x"00", -- $0ddc9
          56778 => x"00", -- $0ddca
          56779 => x"00", -- $0ddcb
          56780 => x"00", -- $0ddcc
          56781 => x"00", -- $0ddcd
          56782 => x"00", -- $0ddce
          56783 => x"00", -- $0ddcf
          56784 => x"00", -- $0ddd0
          56785 => x"00", -- $0ddd1
          56786 => x"00", -- $0ddd2
          56787 => x"00", -- $0ddd3
          56788 => x"00", -- $0ddd4
          56789 => x"00", -- $0ddd5
          56790 => x"00", -- $0ddd6
          56791 => x"00", -- $0ddd7
          56792 => x"00", -- $0ddd8
          56793 => x"00", -- $0ddd9
          56794 => x"00", -- $0ddda
          56795 => x"00", -- $0dddb
          56796 => x"00", -- $0dddc
          56797 => x"00", -- $0dddd
          56798 => x"00", -- $0ddde
          56799 => x"00", -- $0dddf
          56800 => x"00", -- $0dde0
          56801 => x"00", -- $0dde1
          56802 => x"00", -- $0dde2
          56803 => x"00", -- $0dde3
          56804 => x"00", -- $0dde4
          56805 => x"00", -- $0dde5
          56806 => x"00", -- $0dde6
          56807 => x"00", -- $0dde7
          56808 => x"00", -- $0dde8
          56809 => x"00", -- $0dde9
          56810 => x"00", -- $0ddea
          56811 => x"00", -- $0ddeb
          56812 => x"00", -- $0ddec
          56813 => x"00", -- $0dded
          56814 => x"00", -- $0ddee
          56815 => x"00", -- $0ddef
          56816 => x"00", -- $0ddf0
          56817 => x"00", -- $0ddf1
          56818 => x"00", -- $0ddf2
          56819 => x"00", -- $0ddf3
          56820 => x"00", -- $0ddf4
          56821 => x"00", -- $0ddf5
          56822 => x"00", -- $0ddf6
          56823 => x"00", -- $0ddf7
          56824 => x"00", -- $0ddf8
          56825 => x"00", -- $0ddf9
          56826 => x"00", -- $0ddfa
          56827 => x"00", -- $0ddfb
          56828 => x"00", -- $0ddfc
          56829 => x"00", -- $0ddfd
          56830 => x"00", -- $0ddfe
          56831 => x"00", -- $0ddff
          56832 => x"00", -- $0de00
          56833 => x"00", -- $0de01
          56834 => x"00", -- $0de02
          56835 => x"00", -- $0de03
          56836 => x"00", -- $0de04
          56837 => x"00", -- $0de05
          56838 => x"00", -- $0de06
          56839 => x"00", -- $0de07
          56840 => x"00", -- $0de08
          56841 => x"00", -- $0de09
          56842 => x"00", -- $0de0a
          56843 => x"00", -- $0de0b
          56844 => x"00", -- $0de0c
          56845 => x"00", -- $0de0d
          56846 => x"00", -- $0de0e
          56847 => x"00", -- $0de0f
          56848 => x"00", -- $0de10
          56849 => x"00", -- $0de11
          56850 => x"00", -- $0de12
          56851 => x"00", -- $0de13
          56852 => x"00", -- $0de14
          56853 => x"00", -- $0de15
          56854 => x"00", -- $0de16
          56855 => x"00", -- $0de17
          56856 => x"00", -- $0de18
          56857 => x"00", -- $0de19
          56858 => x"00", -- $0de1a
          56859 => x"00", -- $0de1b
          56860 => x"00", -- $0de1c
          56861 => x"00", -- $0de1d
          56862 => x"00", -- $0de1e
          56863 => x"00", -- $0de1f
          56864 => x"00", -- $0de20
          56865 => x"00", -- $0de21
          56866 => x"00", -- $0de22
          56867 => x"00", -- $0de23
          56868 => x"00", -- $0de24
          56869 => x"00", -- $0de25
          56870 => x"00", -- $0de26
          56871 => x"00", -- $0de27
          56872 => x"00", -- $0de28
          56873 => x"00", -- $0de29
          56874 => x"00", -- $0de2a
          56875 => x"00", -- $0de2b
          56876 => x"00", -- $0de2c
          56877 => x"00", -- $0de2d
          56878 => x"00", -- $0de2e
          56879 => x"00", -- $0de2f
          56880 => x"00", -- $0de30
          56881 => x"00", -- $0de31
          56882 => x"00", -- $0de32
          56883 => x"00", -- $0de33
          56884 => x"00", -- $0de34
          56885 => x"00", -- $0de35
          56886 => x"00", -- $0de36
          56887 => x"00", -- $0de37
          56888 => x"00", -- $0de38
          56889 => x"00", -- $0de39
          56890 => x"00", -- $0de3a
          56891 => x"00", -- $0de3b
          56892 => x"00", -- $0de3c
          56893 => x"00", -- $0de3d
          56894 => x"00", -- $0de3e
          56895 => x"00", -- $0de3f
          56896 => x"00", -- $0de40
          56897 => x"00", -- $0de41
          56898 => x"00", -- $0de42
          56899 => x"00", -- $0de43
          56900 => x"00", -- $0de44
          56901 => x"00", -- $0de45
          56902 => x"00", -- $0de46
          56903 => x"00", -- $0de47
          56904 => x"00", -- $0de48
          56905 => x"00", -- $0de49
          56906 => x"00", -- $0de4a
          56907 => x"00", -- $0de4b
          56908 => x"00", -- $0de4c
          56909 => x"00", -- $0de4d
          56910 => x"00", -- $0de4e
          56911 => x"00", -- $0de4f
          56912 => x"00", -- $0de50
          56913 => x"00", -- $0de51
          56914 => x"00", -- $0de52
          56915 => x"00", -- $0de53
          56916 => x"00", -- $0de54
          56917 => x"00", -- $0de55
          56918 => x"00", -- $0de56
          56919 => x"00", -- $0de57
          56920 => x"00", -- $0de58
          56921 => x"00", -- $0de59
          56922 => x"00", -- $0de5a
          56923 => x"00", -- $0de5b
          56924 => x"00", -- $0de5c
          56925 => x"00", -- $0de5d
          56926 => x"00", -- $0de5e
          56927 => x"00", -- $0de5f
          56928 => x"00", -- $0de60
          56929 => x"00", -- $0de61
          56930 => x"00", -- $0de62
          56931 => x"00", -- $0de63
          56932 => x"00", -- $0de64
          56933 => x"00", -- $0de65
          56934 => x"00", -- $0de66
          56935 => x"00", -- $0de67
          56936 => x"00", -- $0de68
          56937 => x"00", -- $0de69
          56938 => x"00", -- $0de6a
          56939 => x"00", -- $0de6b
          56940 => x"00", -- $0de6c
          56941 => x"00", -- $0de6d
          56942 => x"00", -- $0de6e
          56943 => x"00", -- $0de6f
          56944 => x"00", -- $0de70
          56945 => x"00", -- $0de71
          56946 => x"00", -- $0de72
          56947 => x"00", -- $0de73
          56948 => x"00", -- $0de74
          56949 => x"00", -- $0de75
          56950 => x"00", -- $0de76
          56951 => x"00", -- $0de77
          56952 => x"00", -- $0de78
          56953 => x"00", -- $0de79
          56954 => x"00", -- $0de7a
          56955 => x"00", -- $0de7b
          56956 => x"00", -- $0de7c
          56957 => x"00", -- $0de7d
          56958 => x"00", -- $0de7e
          56959 => x"00", -- $0de7f
          56960 => x"00", -- $0de80
          56961 => x"00", -- $0de81
          56962 => x"00", -- $0de82
          56963 => x"00", -- $0de83
          56964 => x"00", -- $0de84
          56965 => x"00", -- $0de85
          56966 => x"00", -- $0de86
          56967 => x"00", -- $0de87
          56968 => x"00", -- $0de88
          56969 => x"00", -- $0de89
          56970 => x"00", -- $0de8a
          56971 => x"00", -- $0de8b
          56972 => x"00", -- $0de8c
          56973 => x"00", -- $0de8d
          56974 => x"00", -- $0de8e
          56975 => x"00", -- $0de8f
          56976 => x"00", -- $0de90
          56977 => x"00", -- $0de91
          56978 => x"00", -- $0de92
          56979 => x"00", -- $0de93
          56980 => x"00", -- $0de94
          56981 => x"00", -- $0de95
          56982 => x"00", -- $0de96
          56983 => x"00", -- $0de97
          56984 => x"00", -- $0de98
          56985 => x"00", -- $0de99
          56986 => x"00", -- $0de9a
          56987 => x"00", -- $0de9b
          56988 => x"00", -- $0de9c
          56989 => x"00", -- $0de9d
          56990 => x"00", -- $0de9e
          56991 => x"00", -- $0de9f
          56992 => x"00", -- $0dea0
          56993 => x"00", -- $0dea1
          56994 => x"00", -- $0dea2
          56995 => x"00", -- $0dea3
          56996 => x"00", -- $0dea4
          56997 => x"00", -- $0dea5
          56998 => x"00", -- $0dea6
          56999 => x"00", -- $0dea7
          57000 => x"00", -- $0dea8
          57001 => x"00", -- $0dea9
          57002 => x"00", -- $0deaa
          57003 => x"00", -- $0deab
          57004 => x"00", -- $0deac
          57005 => x"00", -- $0dead
          57006 => x"00", -- $0deae
          57007 => x"00", -- $0deaf
          57008 => x"00", -- $0deb0
          57009 => x"00", -- $0deb1
          57010 => x"00", -- $0deb2
          57011 => x"00", -- $0deb3
          57012 => x"00", -- $0deb4
          57013 => x"00", -- $0deb5
          57014 => x"00", -- $0deb6
          57015 => x"00", -- $0deb7
          57016 => x"00", -- $0deb8
          57017 => x"00", -- $0deb9
          57018 => x"00", -- $0deba
          57019 => x"00", -- $0debb
          57020 => x"00", -- $0debc
          57021 => x"00", -- $0debd
          57022 => x"00", -- $0debe
          57023 => x"00", -- $0debf
          57024 => x"00", -- $0dec0
          57025 => x"00", -- $0dec1
          57026 => x"00", -- $0dec2
          57027 => x"00", -- $0dec3
          57028 => x"00", -- $0dec4
          57029 => x"00", -- $0dec5
          57030 => x"00", -- $0dec6
          57031 => x"00", -- $0dec7
          57032 => x"00", -- $0dec8
          57033 => x"00", -- $0dec9
          57034 => x"00", -- $0deca
          57035 => x"00", -- $0decb
          57036 => x"00", -- $0decc
          57037 => x"00", -- $0decd
          57038 => x"00", -- $0dece
          57039 => x"00", -- $0decf
          57040 => x"00", -- $0ded0
          57041 => x"00", -- $0ded1
          57042 => x"00", -- $0ded2
          57043 => x"00", -- $0ded3
          57044 => x"00", -- $0ded4
          57045 => x"00", -- $0ded5
          57046 => x"00", -- $0ded6
          57047 => x"00", -- $0ded7
          57048 => x"00", -- $0ded8
          57049 => x"00", -- $0ded9
          57050 => x"00", -- $0deda
          57051 => x"00", -- $0dedb
          57052 => x"00", -- $0dedc
          57053 => x"00", -- $0dedd
          57054 => x"00", -- $0dede
          57055 => x"00", -- $0dedf
          57056 => x"00", -- $0dee0
          57057 => x"00", -- $0dee1
          57058 => x"00", -- $0dee2
          57059 => x"00", -- $0dee3
          57060 => x"00", -- $0dee4
          57061 => x"00", -- $0dee5
          57062 => x"00", -- $0dee6
          57063 => x"00", -- $0dee7
          57064 => x"00", -- $0dee8
          57065 => x"00", -- $0dee9
          57066 => x"00", -- $0deea
          57067 => x"00", -- $0deeb
          57068 => x"00", -- $0deec
          57069 => x"00", -- $0deed
          57070 => x"00", -- $0deee
          57071 => x"00", -- $0deef
          57072 => x"00", -- $0def0
          57073 => x"00", -- $0def1
          57074 => x"00", -- $0def2
          57075 => x"00", -- $0def3
          57076 => x"00", -- $0def4
          57077 => x"00", -- $0def5
          57078 => x"00", -- $0def6
          57079 => x"00", -- $0def7
          57080 => x"00", -- $0def8
          57081 => x"00", -- $0def9
          57082 => x"00", -- $0defa
          57083 => x"00", -- $0defb
          57084 => x"00", -- $0defc
          57085 => x"00", -- $0defd
          57086 => x"00", -- $0defe
          57087 => x"00", -- $0deff
          57088 => x"00", -- $0df00
          57089 => x"00", -- $0df01
          57090 => x"00", -- $0df02
          57091 => x"00", -- $0df03
          57092 => x"00", -- $0df04
          57093 => x"00", -- $0df05
          57094 => x"00", -- $0df06
          57095 => x"00", -- $0df07
          57096 => x"00", -- $0df08
          57097 => x"00", -- $0df09
          57098 => x"00", -- $0df0a
          57099 => x"00", -- $0df0b
          57100 => x"00", -- $0df0c
          57101 => x"00", -- $0df0d
          57102 => x"00", -- $0df0e
          57103 => x"00", -- $0df0f
          57104 => x"00", -- $0df10
          57105 => x"00", -- $0df11
          57106 => x"00", -- $0df12
          57107 => x"00", -- $0df13
          57108 => x"00", -- $0df14
          57109 => x"00", -- $0df15
          57110 => x"00", -- $0df16
          57111 => x"00", -- $0df17
          57112 => x"00", -- $0df18
          57113 => x"00", -- $0df19
          57114 => x"00", -- $0df1a
          57115 => x"00", -- $0df1b
          57116 => x"00", -- $0df1c
          57117 => x"00", -- $0df1d
          57118 => x"00", -- $0df1e
          57119 => x"00", -- $0df1f
          57120 => x"00", -- $0df20
          57121 => x"00", -- $0df21
          57122 => x"00", -- $0df22
          57123 => x"00", -- $0df23
          57124 => x"00", -- $0df24
          57125 => x"00", -- $0df25
          57126 => x"00", -- $0df26
          57127 => x"00", -- $0df27
          57128 => x"00", -- $0df28
          57129 => x"00", -- $0df29
          57130 => x"00", -- $0df2a
          57131 => x"00", -- $0df2b
          57132 => x"00", -- $0df2c
          57133 => x"00", -- $0df2d
          57134 => x"00", -- $0df2e
          57135 => x"00", -- $0df2f
          57136 => x"00", -- $0df30
          57137 => x"00", -- $0df31
          57138 => x"00", -- $0df32
          57139 => x"00", -- $0df33
          57140 => x"00", -- $0df34
          57141 => x"00", -- $0df35
          57142 => x"00", -- $0df36
          57143 => x"00", -- $0df37
          57144 => x"00", -- $0df38
          57145 => x"00", -- $0df39
          57146 => x"00", -- $0df3a
          57147 => x"00", -- $0df3b
          57148 => x"00", -- $0df3c
          57149 => x"00", -- $0df3d
          57150 => x"00", -- $0df3e
          57151 => x"00", -- $0df3f
          57152 => x"00", -- $0df40
          57153 => x"00", -- $0df41
          57154 => x"00", -- $0df42
          57155 => x"00", -- $0df43
          57156 => x"00", -- $0df44
          57157 => x"00", -- $0df45
          57158 => x"00", -- $0df46
          57159 => x"00", -- $0df47
          57160 => x"00", -- $0df48
          57161 => x"00", -- $0df49
          57162 => x"00", -- $0df4a
          57163 => x"00", -- $0df4b
          57164 => x"00", -- $0df4c
          57165 => x"00", -- $0df4d
          57166 => x"00", -- $0df4e
          57167 => x"00", -- $0df4f
          57168 => x"00", -- $0df50
          57169 => x"00", -- $0df51
          57170 => x"00", -- $0df52
          57171 => x"00", -- $0df53
          57172 => x"00", -- $0df54
          57173 => x"00", -- $0df55
          57174 => x"00", -- $0df56
          57175 => x"00", -- $0df57
          57176 => x"00", -- $0df58
          57177 => x"00", -- $0df59
          57178 => x"00", -- $0df5a
          57179 => x"00", -- $0df5b
          57180 => x"00", -- $0df5c
          57181 => x"00", -- $0df5d
          57182 => x"00", -- $0df5e
          57183 => x"00", -- $0df5f
          57184 => x"00", -- $0df60
          57185 => x"00", -- $0df61
          57186 => x"00", -- $0df62
          57187 => x"00", -- $0df63
          57188 => x"00", -- $0df64
          57189 => x"00", -- $0df65
          57190 => x"00", -- $0df66
          57191 => x"00", -- $0df67
          57192 => x"00", -- $0df68
          57193 => x"00", -- $0df69
          57194 => x"00", -- $0df6a
          57195 => x"00", -- $0df6b
          57196 => x"00", -- $0df6c
          57197 => x"00", -- $0df6d
          57198 => x"00", -- $0df6e
          57199 => x"00", -- $0df6f
          57200 => x"00", -- $0df70
          57201 => x"00", -- $0df71
          57202 => x"00", -- $0df72
          57203 => x"00", -- $0df73
          57204 => x"00", -- $0df74
          57205 => x"00", -- $0df75
          57206 => x"00", -- $0df76
          57207 => x"00", -- $0df77
          57208 => x"00", -- $0df78
          57209 => x"00", -- $0df79
          57210 => x"00", -- $0df7a
          57211 => x"00", -- $0df7b
          57212 => x"00", -- $0df7c
          57213 => x"00", -- $0df7d
          57214 => x"00", -- $0df7e
          57215 => x"00", -- $0df7f
          57216 => x"00", -- $0df80
          57217 => x"00", -- $0df81
          57218 => x"00", -- $0df82
          57219 => x"00", -- $0df83
          57220 => x"00", -- $0df84
          57221 => x"00", -- $0df85
          57222 => x"00", -- $0df86
          57223 => x"00", -- $0df87
          57224 => x"00", -- $0df88
          57225 => x"00", -- $0df89
          57226 => x"00", -- $0df8a
          57227 => x"00", -- $0df8b
          57228 => x"00", -- $0df8c
          57229 => x"00", -- $0df8d
          57230 => x"00", -- $0df8e
          57231 => x"00", -- $0df8f
          57232 => x"00", -- $0df90
          57233 => x"00", -- $0df91
          57234 => x"00", -- $0df92
          57235 => x"00", -- $0df93
          57236 => x"00", -- $0df94
          57237 => x"00", -- $0df95
          57238 => x"00", -- $0df96
          57239 => x"00", -- $0df97
          57240 => x"00", -- $0df98
          57241 => x"00", -- $0df99
          57242 => x"00", -- $0df9a
          57243 => x"00", -- $0df9b
          57244 => x"00", -- $0df9c
          57245 => x"00", -- $0df9d
          57246 => x"00", -- $0df9e
          57247 => x"00", -- $0df9f
          57248 => x"00", -- $0dfa0
          57249 => x"00", -- $0dfa1
          57250 => x"00", -- $0dfa2
          57251 => x"00", -- $0dfa3
          57252 => x"00", -- $0dfa4
          57253 => x"00", -- $0dfa5
          57254 => x"00", -- $0dfa6
          57255 => x"00", -- $0dfa7
          57256 => x"00", -- $0dfa8
          57257 => x"00", -- $0dfa9
          57258 => x"00", -- $0dfaa
          57259 => x"00", -- $0dfab
          57260 => x"00", -- $0dfac
          57261 => x"00", -- $0dfad
          57262 => x"00", -- $0dfae
          57263 => x"00", -- $0dfaf
          57264 => x"00", -- $0dfb0
          57265 => x"00", -- $0dfb1
          57266 => x"00", -- $0dfb2
          57267 => x"00", -- $0dfb3
          57268 => x"00", -- $0dfb4
          57269 => x"00", -- $0dfb5
          57270 => x"00", -- $0dfb6
          57271 => x"00", -- $0dfb7
          57272 => x"00", -- $0dfb8
          57273 => x"00", -- $0dfb9
          57274 => x"00", -- $0dfba
          57275 => x"00", -- $0dfbb
          57276 => x"00", -- $0dfbc
          57277 => x"00", -- $0dfbd
          57278 => x"00", -- $0dfbe
          57279 => x"00", -- $0dfbf
          57280 => x"00", -- $0dfc0
          57281 => x"00", -- $0dfc1
          57282 => x"00", -- $0dfc2
          57283 => x"00", -- $0dfc3
          57284 => x"00", -- $0dfc4
          57285 => x"00", -- $0dfc5
          57286 => x"00", -- $0dfc6
          57287 => x"00", -- $0dfc7
          57288 => x"00", -- $0dfc8
          57289 => x"00", -- $0dfc9
          57290 => x"00", -- $0dfca
          57291 => x"00", -- $0dfcb
          57292 => x"00", -- $0dfcc
          57293 => x"00", -- $0dfcd
          57294 => x"00", -- $0dfce
          57295 => x"00", -- $0dfcf
          57296 => x"00", -- $0dfd0
          57297 => x"00", -- $0dfd1
          57298 => x"00", -- $0dfd2
          57299 => x"00", -- $0dfd3
          57300 => x"00", -- $0dfd4
          57301 => x"00", -- $0dfd5
          57302 => x"00", -- $0dfd6
          57303 => x"00", -- $0dfd7
          57304 => x"00", -- $0dfd8
          57305 => x"00", -- $0dfd9
          57306 => x"00", -- $0dfda
          57307 => x"00", -- $0dfdb
          57308 => x"00", -- $0dfdc
          57309 => x"00", -- $0dfdd
          57310 => x"00", -- $0dfde
          57311 => x"00", -- $0dfdf
          57312 => x"00", -- $0dfe0
          57313 => x"00", -- $0dfe1
          57314 => x"00", -- $0dfe2
          57315 => x"00", -- $0dfe3
          57316 => x"00", -- $0dfe4
          57317 => x"00", -- $0dfe5
          57318 => x"00", -- $0dfe6
          57319 => x"00", -- $0dfe7
          57320 => x"00", -- $0dfe8
          57321 => x"00", -- $0dfe9
          57322 => x"00", -- $0dfea
          57323 => x"00", -- $0dfeb
          57324 => x"00", -- $0dfec
          57325 => x"00", -- $0dfed
          57326 => x"00", -- $0dfee
          57327 => x"00", -- $0dfef
          57328 => x"00", -- $0dff0
          57329 => x"00", -- $0dff1
          57330 => x"00", -- $0dff2
          57331 => x"00", -- $0dff3
          57332 => x"00", -- $0dff4
          57333 => x"00", -- $0dff5
          57334 => x"00", -- $0dff6
          57335 => x"00", -- $0dff7
          57336 => x"00", -- $0dff8
          57337 => x"00", -- $0dff9
          57338 => x"00", -- $0dffa
          57339 => x"00", -- $0dffb
          57340 => x"00", -- $0dffc
          57341 => x"00", -- $0dffd
          57342 => x"00", -- $0dffe
          57343 => x"00", -- $0dfff
          57344 => x"00", -- $0e000
          57345 => x"00", -- $0e001
          57346 => x"00", -- $0e002
          57347 => x"00", -- $0e003
          57348 => x"00", -- $0e004
          57349 => x"00", -- $0e005
          57350 => x"00", -- $0e006
          57351 => x"00", -- $0e007
          57352 => x"00", -- $0e008
          57353 => x"00", -- $0e009
          57354 => x"00", -- $0e00a
          57355 => x"00", -- $0e00b
          57356 => x"00", -- $0e00c
          57357 => x"00", -- $0e00d
          57358 => x"00", -- $0e00e
          57359 => x"00", -- $0e00f
          57360 => x"00", -- $0e010
          57361 => x"00", -- $0e011
          57362 => x"00", -- $0e012
          57363 => x"00", -- $0e013
          57364 => x"00", -- $0e014
          57365 => x"00", -- $0e015
          57366 => x"00", -- $0e016
          57367 => x"00", -- $0e017
          57368 => x"00", -- $0e018
          57369 => x"00", -- $0e019
          57370 => x"00", -- $0e01a
          57371 => x"00", -- $0e01b
          57372 => x"00", -- $0e01c
          57373 => x"00", -- $0e01d
          57374 => x"00", -- $0e01e
          57375 => x"00", -- $0e01f
          57376 => x"00", -- $0e020
          57377 => x"00", -- $0e021
          57378 => x"00", -- $0e022
          57379 => x"00", -- $0e023
          57380 => x"00", -- $0e024
          57381 => x"00", -- $0e025
          57382 => x"00", -- $0e026
          57383 => x"00", -- $0e027
          57384 => x"00", -- $0e028
          57385 => x"00", -- $0e029
          57386 => x"00", -- $0e02a
          57387 => x"00", -- $0e02b
          57388 => x"00", -- $0e02c
          57389 => x"00", -- $0e02d
          57390 => x"00", -- $0e02e
          57391 => x"00", -- $0e02f
          57392 => x"00", -- $0e030
          57393 => x"00", -- $0e031
          57394 => x"00", -- $0e032
          57395 => x"00", -- $0e033
          57396 => x"00", -- $0e034
          57397 => x"00", -- $0e035
          57398 => x"00", -- $0e036
          57399 => x"00", -- $0e037
          57400 => x"00", -- $0e038
          57401 => x"00", -- $0e039
          57402 => x"00", -- $0e03a
          57403 => x"00", -- $0e03b
          57404 => x"00", -- $0e03c
          57405 => x"00", -- $0e03d
          57406 => x"00", -- $0e03e
          57407 => x"00", -- $0e03f
          57408 => x"00", -- $0e040
          57409 => x"00", -- $0e041
          57410 => x"00", -- $0e042
          57411 => x"00", -- $0e043
          57412 => x"00", -- $0e044
          57413 => x"00", -- $0e045
          57414 => x"00", -- $0e046
          57415 => x"00", -- $0e047
          57416 => x"00", -- $0e048
          57417 => x"00", -- $0e049
          57418 => x"00", -- $0e04a
          57419 => x"00", -- $0e04b
          57420 => x"00", -- $0e04c
          57421 => x"00", -- $0e04d
          57422 => x"00", -- $0e04e
          57423 => x"00", -- $0e04f
          57424 => x"00", -- $0e050
          57425 => x"00", -- $0e051
          57426 => x"00", -- $0e052
          57427 => x"00", -- $0e053
          57428 => x"00", -- $0e054
          57429 => x"00", -- $0e055
          57430 => x"00", -- $0e056
          57431 => x"00", -- $0e057
          57432 => x"00", -- $0e058
          57433 => x"00", -- $0e059
          57434 => x"00", -- $0e05a
          57435 => x"00", -- $0e05b
          57436 => x"00", -- $0e05c
          57437 => x"00", -- $0e05d
          57438 => x"00", -- $0e05e
          57439 => x"00", -- $0e05f
          57440 => x"00", -- $0e060
          57441 => x"00", -- $0e061
          57442 => x"00", -- $0e062
          57443 => x"00", -- $0e063
          57444 => x"00", -- $0e064
          57445 => x"00", -- $0e065
          57446 => x"00", -- $0e066
          57447 => x"00", -- $0e067
          57448 => x"00", -- $0e068
          57449 => x"00", -- $0e069
          57450 => x"00", -- $0e06a
          57451 => x"00", -- $0e06b
          57452 => x"00", -- $0e06c
          57453 => x"00", -- $0e06d
          57454 => x"00", -- $0e06e
          57455 => x"00", -- $0e06f
          57456 => x"00", -- $0e070
          57457 => x"00", -- $0e071
          57458 => x"00", -- $0e072
          57459 => x"00", -- $0e073
          57460 => x"00", -- $0e074
          57461 => x"00", -- $0e075
          57462 => x"00", -- $0e076
          57463 => x"00", -- $0e077
          57464 => x"00", -- $0e078
          57465 => x"00", -- $0e079
          57466 => x"00", -- $0e07a
          57467 => x"00", -- $0e07b
          57468 => x"00", -- $0e07c
          57469 => x"00", -- $0e07d
          57470 => x"00", -- $0e07e
          57471 => x"00", -- $0e07f
          57472 => x"00", -- $0e080
          57473 => x"00", -- $0e081
          57474 => x"00", -- $0e082
          57475 => x"00", -- $0e083
          57476 => x"00", -- $0e084
          57477 => x"00", -- $0e085
          57478 => x"00", -- $0e086
          57479 => x"00", -- $0e087
          57480 => x"00", -- $0e088
          57481 => x"00", -- $0e089
          57482 => x"00", -- $0e08a
          57483 => x"00", -- $0e08b
          57484 => x"00", -- $0e08c
          57485 => x"00", -- $0e08d
          57486 => x"00", -- $0e08e
          57487 => x"00", -- $0e08f
          57488 => x"00", -- $0e090
          57489 => x"00", -- $0e091
          57490 => x"00", -- $0e092
          57491 => x"00", -- $0e093
          57492 => x"00", -- $0e094
          57493 => x"00", -- $0e095
          57494 => x"00", -- $0e096
          57495 => x"00", -- $0e097
          57496 => x"00", -- $0e098
          57497 => x"00", -- $0e099
          57498 => x"00", -- $0e09a
          57499 => x"00", -- $0e09b
          57500 => x"00", -- $0e09c
          57501 => x"00", -- $0e09d
          57502 => x"00", -- $0e09e
          57503 => x"00", -- $0e09f
          57504 => x"00", -- $0e0a0
          57505 => x"00", -- $0e0a1
          57506 => x"00", -- $0e0a2
          57507 => x"00", -- $0e0a3
          57508 => x"00", -- $0e0a4
          57509 => x"00", -- $0e0a5
          57510 => x"00", -- $0e0a6
          57511 => x"00", -- $0e0a7
          57512 => x"00", -- $0e0a8
          57513 => x"00", -- $0e0a9
          57514 => x"00", -- $0e0aa
          57515 => x"00", -- $0e0ab
          57516 => x"00", -- $0e0ac
          57517 => x"00", -- $0e0ad
          57518 => x"00", -- $0e0ae
          57519 => x"00", -- $0e0af
          57520 => x"00", -- $0e0b0
          57521 => x"00", -- $0e0b1
          57522 => x"00", -- $0e0b2
          57523 => x"00", -- $0e0b3
          57524 => x"00", -- $0e0b4
          57525 => x"00", -- $0e0b5
          57526 => x"00", -- $0e0b6
          57527 => x"00", -- $0e0b7
          57528 => x"00", -- $0e0b8
          57529 => x"00", -- $0e0b9
          57530 => x"00", -- $0e0ba
          57531 => x"00", -- $0e0bb
          57532 => x"00", -- $0e0bc
          57533 => x"00", -- $0e0bd
          57534 => x"00", -- $0e0be
          57535 => x"00", -- $0e0bf
          57536 => x"00", -- $0e0c0
          57537 => x"00", -- $0e0c1
          57538 => x"00", -- $0e0c2
          57539 => x"00", -- $0e0c3
          57540 => x"00", -- $0e0c4
          57541 => x"00", -- $0e0c5
          57542 => x"00", -- $0e0c6
          57543 => x"00", -- $0e0c7
          57544 => x"00", -- $0e0c8
          57545 => x"00", -- $0e0c9
          57546 => x"00", -- $0e0ca
          57547 => x"00", -- $0e0cb
          57548 => x"00", -- $0e0cc
          57549 => x"00", -- $0e0cd
          57550 => x"00", -- $0e0ce
          57551 => x"00", -- $0e0cf
          57552 => x"00", -- $0e0d0
          57553 => x"00", -- $0e0d1
          57554 => x"00", -- $0e0d2
          57555 => x"00", -- $0e0d3
          57556 => x"00", -- $0e0d4
          57557 => x"00", -- $0e0d5
          57558 => x"00", -- $0e0d6
          57559 => x"00", -- $0e0d7
          57560 => x"00", -- $0e0d8
          57561 => x"00", -- $0e0d9
          57562 => x"00", -- $0e0da
          57563 => x"00", -- $0e0db
          57564 => x"00", -- $0e0dc
          57565 => x"00", -- $0e0dd
          57566 => x"00", -- $0e0de
          57567 => x"00", -- $0e0df
          57568 => x"00", -- $0e0e0
          57569 => x"00", -- $0e0e1
          57570 => x"00", -- $0e0e2
          57571 => x"00", -- $0e0e3
          57572 => x"00", -- $0e0e4
          57573 => x"00", -- $0e0e5
          57574 => x"00", -- $0e0e6
          57575 => x"00", -- $0e0e7
          57576 => x"00", -- $0e0e8
          57577 => x"00", -- $0e0e9
          57578 => x"00", -- $0e0ea
          57579 => x"00", -- $0e0eb
          57580 => x"00", -- $0e0ec
          57581 => x"00", -- $0e0ed
          57582 => x"00", -- $0e0ee
          57583 => x"00", -- $0e0ef
          57584 => x"00", -- $0e0f0
          57585 => x"00", -- $0e0f1
          57586 => x"00", -- $0e0f2
          57587 => x"00", -- $0e0f3
          57588 => x"00", -- $0e0f4
          57589 => x"00", -- $0e0f5
          57590 => x"00", -- $0e0f6
          57591 => x"00", -- $0e0f7
          57592 => x"00", -- $0e0f8
          57593 => x"00", -- $0e0f9
          57594 => x"00", -- $0e0fa
          57595 => x"00", -- $0e0fb
          57596 => x"00", -- $0e0fc
          57597 => x"00", -- $0e0fd
          57598 => x"00", -- $0e0fe
          57599 => x"00", -- $0e0ff
          57600 => x"00", -- $0e100
          57601 => x"00", -- $0e101
          57602 => x"00", -- $0e102
          57603 => x"00", -- $0e103
          57604 => x"00", -- $0e104
          57605 => x"00", -- $0e105
          57606 => x"00", -- $0e106
          57607 => x"00", -- $0e107
          57608 => x"00", -- $0e108
          57609 => x"00", -- $0e109
          57610 => x"00", -- $0e10a
          57611 => x"00", -- $0e10b
          57612 => x"00", -- $0e10c
          57613 => x"00", -- $0e10d
          57614 => x"00", -- $0e10e
          57615 => x"00", -- $0e10f
          57616 => x"00", -- $0e110
          57617 => x"00", -- $0e111
          57618 => x"00", -- $0e112
          57619 => x"00", -- $0e113
          57620 => x"00", -- $0e114
          57621 => x"00", -- $0e115
          57622 => x"00", -- $0e116
          57623 => x"00", -- $0e117
          57624 => x"00", -- $0e118
          57625 => x"00", -- $0e119
          57626 => x"00", -- $0e11a
          57627 => x"00", -- $0e11b
          57628 => x"00", -- $0e11c
          57629 => x"00", -- $0e11d
          57630 => x"00", -- $0e11e
          57631 => x"00", -- $0e11f
          57632 => x"00", -- $0e120
          57633 => x"00", -- $0e121
          57634 => x"00", -- $0e122
          57635 => x"00", -- $0e123
          57636 => x"00", -- $0e124
          57637 => x"00", -- $0e125
          57638 => x"00", -- $0e126
          57639 => x"00", -- $0e127
          57640 => x"00", -- $0e128
          57641 => x"00", -- $0e129
          57642 => x"00", -- $0e12a
          57643 => x"00", -- $0e12b
          57644 => x"00", -- $0e12c
          57645 => x"00", -- $0e12d
          57646 => x"00", -- $0e12e
          57647 => x"00", -- $0e12f
          57648 => x"00", -- $0e130
          57649 => x"00", -- $0e131
          57650 => x"00", -- $0e132
          57651 => x"00", -- $0e133
          57652 => x"00", -- $0e134
          57653 => x"00", -- $0e135
          57654 => x"00", -- $0e136
          57655 => x"00", -- $0e137
          57656 => x"00", -- $0e138
          57657 => x"00", -- $0e139
          57658 => x"00", -- $0e13a
          57659 => x"00", -- $0e13b
          57660 => x"00", -- $0e13c
          57661 => x"00", -- $0e13d
          57662 => x"00", -- $0e13e
          57663 => x"00", -- $0e13f
          57664 => x"00", -- $0e140
          57665 => x"00", -- $0e141
          57666 => x"00", -- $0e142
          57667 => x"00", -- $0e143
          57668 => x"00", -- $0e144
          57669 => x"00", -- $0e145
          57670 => x"00", -- $0e146
          57671 => x"00", -- $0e147
          57672 => x"00", -- $0e148
          57673 => x"00", -- $0e149
          57674 => x"00", -- $0e14a
          57675 => x"00", -- $0e14b
          57676 => x"00", -- $0e14c
          57677 => x"00", -- $0e14d
          57678 => x"00", -- $0e14e
          57679 => x"00", -- $0e14f
          57680 => x"00", -- $0e150
          57681 => x"00", -- $0e151
          57682 => x"00", -- $0e152
          57683 => x"00", -- $0e153
          57684 => x"00", -- $0e154
          57685 => x"00", -- $0e155
          57686 => x"00", -- $0e156
          57687 => x"00", -- $0e157
          57688 => x"00", -- $0e158
          57689 => x"00", -- $0e159
          57690 => x"00", -- $0e15a
          57691 => x"00", -- $0e15b
          57692 => x"00", -- $0e15c
          57693 => x"00", -- $0e15d
          57694 => x"00", -- $0e15e
          57695 => x"00", -- $0e15f
          57696 => x"00", -- $0e160
          57697 => x"00", -- $0e161
          57698 => x"00", -- $0e162
          57699 => x"00", -- $0e163
          57700 => x"00", -- $0e164
          57701 => x"00", -- $0e165
          57702 => x"00", -- $0e166
          57703 => x"00", -- $0e167
          57704 => x"00", -- $0e168
          57705 => x"00", -- $0e169
          57706 => x"00", -- $0e16a
          57707 => x"00", -- $0e16b
          57708 => x"00", -- $0e16c
          57709 => x"00", -- $0e16d
          57710 => x"00", -- $0e16e
          57711 => x"00", -- $0e16f
          57712 => x"00", -- $0e170
          57713 => x"00", -- $0e171
          57714 => x"00", -- $0e172
          57715 => x"00", -- $0e173
          57716 => x"00", -- $0e174
          57717 => x"00", -- $0e175
          57718 => x"00", -- $0e176
          57719 => x"00", -- $0e177
          57720 => x"00", -- $0e178
          57721 => x"00", -- $0e179
          57722 => x"00", -- $0e17a
          57723 => x"00", -- $0e17b
          57724 => x"00", -- $0e17c
          57725 => x"00", -- $0e17d
          57726 => x"00", -- $0e17e
          57727 => x"00", -- $0e17f
          57728 => x"00", -- $0e180
          57729 => x"00", -- $0e181
          57730 => x"00", -- $0e182
          57731 => x"00", -- $0e183
          57732 => x"00", -- $0e184
          57733 => x"00", -- $0e185
          57734 => x"00", -- $0e186
          57735 => x"00", -- $0e187
          57736 => x"00", -- $0e188
          57737 => x"00", -- $0e189
          57738 => x"00", -- $0e18a
          57739 => x"00", -- $0e18b
          57740 => x"00", -- $0e18c
          57741 => x"00", -- $0e18d
          57742 => x"00", -- $0e18e
          57743 => x"00", -- $0e18f
          57744 => x"00", -- $0e190
          57745 => x"00", -- $0e191
          57746 => x"00", -- $0e192
          57747 => x"00", -- $0e193
          57748 => x"00", -- $0e194
          57749 => x"00", -- $0e195
          57750 => x"00", -- $0e196
          57751 => x"00", -- $0e197
          57752 => x"00", -- $0e198
          57753 => x"00", -- $0e199
          57754 => x"00", -- $0e19a
          57755 => x"00", -- $0e19b
          57756 => x"00", -- $0e19c
          57757 => x"00", -- $0e19d
          57758 => x"00", -- $0e19e
          57759 => x"00", -- $0e19f
          57760 => x"00", -- $0e1a0
          57761 => x"00", -- $0e1a1
          57762 => x"00", -- $0e1a2
          57763 => x"00", -- $0e1a3
          57764 => x"00", -- $0e1a4
          57765 => x"00", -- $0e1a5
          57766 => x"00", -- $0e1a6
          57767 => x"00", -- $0e1a7
          57768 => x"00", -- $0e1a8
          57769 => x"00", -- $0e1a9
          57770 => x"00", -- $0e1aa
          57771 => x"00", -- $0e1ab
          57772 => x"00", -- $0e1ac
          57773 => x"00", -- $0e1ad
          57774 => x"00", -- $0e1ae
          57775 => x"00", -- $0e1af
          57776 => x"00", -- $0e1b0
          57777 => x"00", -- $0e1b1
          57778 => x"00", -- $0e1b2
          57779 => x"00", -- $0e1b3
          57780 => x"00", -- $0e1b4
          57781 => x"00", -- $0e1b5
          57782 => x"00", -- $0e1b6
          57783 => x"00", -- $0e1b7
          57784 => x"00", -- $0e1b8
          57785 => x"00", -- $0e1b9
          57786 => x"00", -- $0e1ba
          57787 => x"00", -- $0e1bb
          57788 => x"00", -- $0e1bc
          57789 => x"00", -- $0e1bd
          57790 => x"00", -- $0e1be
          57791 => x"00", -- $0e1bf
          57792 => x"00", -- $0e1c0
          57793 => x"00", -- $0e1c1
          57794 => x"00", -- $0e1c2
          57795 => x"00", -- $0e1c3
          57796 => x"00", -- $0e1c4
          57797 => x"00", -- $0e1c5
          57798 => x"00", -- $0e1c6
          57799 => x"00", -- $0e1c7
          57800 => x"00", -- $0e1c8
          57801 => x"00", -- $0e1c9
          57802 => x"00", -- $0e1ca
          57803 => x"00", -- $0e1cb
          57804 => x"00", -- $0e1cc
          57805 => x"00", -- $0e1cd
          57806 => x"00", -- $0e1ce
          57807 => x"00", -- $0e1cf
          57808 => x"00", -- $0e1d0
          57809 => x"00", -- $0e1d1
          57810 => x"00", -- $0e1d2
          57811 => x"00", -- $0e1d3
          57812 => x"00", -- $0e1d4
          57813 => x"00", -- $0e1d5
          57814 => x"00", -- $0e1d6
          57815 => x"00", -- $0e1d7
          57816 => x"00", -- $0e1d8
          57817 => x"00", -- $0e1d9
          57818 => x"00", -- $0e1da
          57819 => x"00", -- $0e1db
          57820 => x"00", -- $0e1dc
          57821 => x"00", -- $0e1dd
          57822 => x"00", -- $0e1de
          57823 => x"00", -- $0e1df
          57824 => x"00", -- $0e1e0
          57825 => x"00", -- $0e1e1
          57826 => x"00", -- $0e1e2
          57827 => x"00", -- $0e1e3
          57828 => x"00", -- $0e1e4
          57829 => x"00", -- $0e1e5
          57830 => x"00", -- $0e1e6
          57831 => x"00", -- $0e1e7
          57832 => x"00", -- $0e1e8
          57833 => x"00", -- $0e1e9
          57834 => x"00", -- $0e1ea
          57835 => x"00", -- $0e1eb
          57836 => x"00", -- $0e1ec
          57837 => x"00", -- $0e1ed
          57838 => x"00", -- $0e1ee
          57839 => x"00", -- $0e1ef
          57840 => x"00", -- $0e1f0
          57841 => x"00", -- $0e1f1
          57842 => x"00", -- $0e1f2
          57843 => x"00", -- $0e1f3
          57844 => x"00", -- $0e1f4
          57845 => x"00", -- $0e1f5
          57846 => x"00", -- $0e1f6
          57847 => x"00", -- $0e1f7
          57848 => x"00", -- $0e1f8
          57849 => x"00", -- $0e1f9
          57850 => x"00", -- $0e1fa
          57851 => x"00", -- $0e1fb
          57852 => x"00", -- $0e1fc
          57853 => x"00", -- $0e1fd
          57854 => x"00", -- $0e1fe
          57855 => x"00", -- $0e1ff
          57856 => x"00", -- $0e200
          57857 => x"00", -- $0e201
          57858 => x"00", -- $0e202
          57859 => x"00", -- $0e203
          57860 => x"00", -- $0e204
          57861 => x"00", -- $0e205
          57862 => x"00", -- $0e206
          57863 => x"00", -- $0e207
          57864 => x"00", -- $0e208
          57865 => x"00", -- $0e209
          57866 => x"00", -- $0e20a
          57867 => x"00", -- $0e20b
          57868 => x"00", -- $0e20c
          57869 => x"00", -- $0e20d
          57870 => x"00", -- $0e20e
          57871 => x"00", -- $0e20f
          57872 => x"00", -- $0e210
          57873 => x"00", -- $0e211
          57874 => x"00", -- $0e212
          57875 => x"00", -- $0e213
          57876 => x"00", -- $0e214
          57877 => x"00", -- $0e215
          57878 => x"00", -- $0e216
          57879 => x"00", -- $0e217
          57880 => x"00", -- $0e218
          57881 => x"00", -- $0e219
          57882 => x"00", -- $0e21a
          57883 => x"00", -- $0e21b
          57884 => x"00", -- $0e21c
          57885 => x"00", -- $0e21d
          57886 => x"00", -- $0e21e
          57887 => x"00", -- $0e21f
          57888 => x"00", -- $0e220
          57889 => x"00", -- $0e221
          57890 => x"00", -- $0e222
          57891 => x"00", -- $0e223
          57892 => x"00", -- $0e224
          57893 => x"00", -- $0e225
          57894 => x"00", -- $0e226
          57895 => x"00", -- $0e227
          57896 => x"00", -- $0e228
          57897 => x"00", -- $0e229
          57898 => x"00", -- $0e22a
          57899 => x"00", -- $0e22b
          57900 => x"00", -- $0e22c
          57901 => x"00", -- $0e22d
          57902 => x"00", -- $0e22e
          57903 => x"00", -- $0e22f
          57904 => x"00", -- $0e230
          57905 => x"00", -- $0e231
          57906 => x"00", -- $0e232
          57907 => x"00", -- $0e233
          57908 => x"00", -- $0e234
          57909 => x"00", -- $0e235
          57910 => x"00", -- $0e236
          57911 => x"00", -- $0e237
          57912 => x"00", -- $0e238
          57913 => x"00", -- $0e239
          57914 => x"00", -- $0e23a
          57915 => x"00", -- $0e23b
          57916 => x"00", -- $0e23c
          57917 => x"00", -- $0e23d
          57918 => x"00", -- $0e23e
          57919 => x"00", -- $0e23f
          57920 => x"00", -- $0e240
          57921 => x"00", -- $0e241
          57922 => x"00", -- $0e242
          57923 => x"00", -- $0e243
          57924 => x"00", -- $0e244
          57925 => x"00", -- $0e245
          57926 => x"00", -- $0e246
          57927 => x"00", -- $0e247
          57928 => x"00", -- $0e248
          57929 => x"00", -- $0e249
          57930 => x"00", -- $0e24a
          57931 => x"00", -- $0e24b
          57932 => x"00", -- $0e24c
          57933 => x"00", -- $0e24d
          57934 => x"00", -- $0e24e
          57935 => x"00", -- $0e24f
          57936 => x"00", -- $0e250
          57937 => x"00", -- $0e251
          57938 => x"00", -- $0e252
          57939 => x"00", -- $0e253
          57940 => x"00", -- $0e254
          57941 => x"00", -- $0e255
          57942 => x"00", -- $0e256
          57943 => x"00", -- $0e257
          57944 => x"00", -- $0e258
          57945 => x"00", -- $0e259
          57946 => x"00", -- $0e25a
          57947 => x"00", -- $0e25b
          57948 => x"00", -- $0e25c
          57949 => x"00", -- $0e25d
          57950 => x"00", -- $0e25e
          57951 => x"00", -- $0e25f
          57952 => x"00", -- $0e260
          57953 => x"00", -- $0e261
          57954 => x"00", -- $0e262
          57955 => x"00", -- $0e263
          57956 => x"00", -- $0e264
          57957 => x"00", -- $0e265
          57958 => x"00", -- $0e266
          57959 => x"00", -- $0e267
          57960 => x"00", -- $0e268
          57961 => x"00", -- $0e269
          57962 => x"00", -- $0e26a
          57963 => x"00", -- $0e26b
          57964 => x"00", -- $0e26c
          57965 => x"00", -- $0e26d
          57966 => x"00", -- $0e26e
          57967 => x"00", -- $0e26f
          57968 => x"00", -- $0e270
          57969 => x"00", -- $0e271
          57970 => x"00", -- $0e272
          57971 => x"00", -- $0e273
          57972 => x"00", -- $0e274
          57973 => x"00", -- $0e275
          57974 => x"00", -- $0e276
          57975 => x"00", -- $0e277
          57976 => x"00", -- $0e278
          57977 => x"00", -- $0e279
          57978 => x"00", -- $0e27a
          57979 => x"00", -- $0e27b
          57980 => x"00", -- $0e27c
          57981 => x"00", -- $0e27d
          57982 => x"00", -- $0e27e
          57983 => x"00", -- $0e27f
          57984 => x"00", -- $0e280
          57985 => x"00", -- $0e281
          57986 => x"00", -- $0e282
          57987 => x"00", -- $0e283
          57988 => x"00", -- $0e284
          57989 => x"00", -- $0e285
          57990 => x"00", -- $0e286
          57991 => x"00", -- $0e287
          57992 => x"00", -- $0e288
          57993 => x"00", -- $0e289
          57994 => x"00", -- $0e28a
          57995 => x"00", -- $0e28b
          57996 => x"00", -- $0e28c
          57997 => x"00", -- $0e28d
          57998 => x"00", -- $0e28e
          57999 => x"00", -- $0e28f
          58000 => x"00", -- $0e290
          58001 => x"00", -- $0e291
          58002 => x"00", -- $0e292
          58003 => x"00", -- $0e293
          58004 => x"00", -- $0e294
          58005 => x"00", -- $0e295
          58006 => x"00", -- $0e296
          58007 => x"00", -- $0e297
          58008 => x"00", -- $0e298
          58009 => x"00", -- $0e299
          58010 => x"00", -- $0e29a
          58011 => x"00", -- $0e29b
          58012 => x"00", -- $0e29c
          58013 => x"00", -- $0e29d
          58014 => x"00", -- $0e29e
          58015 => x"00", -- $0e29f
          58016 => x"00", -- $0e2a0
          58017 => x"00", -- $0e2a1
          58018 => x"00", -- $0e2a2
          58019 => x"00", -- $0e2a3
          58020 => x"00", -- $0e2a4
          58021 => x"00", -- $0e2a5
          58022 => x"00", -- $0e2a6
          58023 => x"00", -- $0e2a7
          58024 => x"00", -- $0e2a8
          58025 => x"00", -- $0e2a9
          58026 => x"00", -- $0e2aa
          58027 => x"00", -- $0e2ab
          58028 => x"00", -- $0e2ac
          58029 => x"00", -- $0e2ad
          58030 => x"00", -- $0e2ae
          58031 => x"00", -- $0e2af
          58032 => x"00", -- $0e2b0
          58033 => x"00", -- $0e2b1
          58034 => x"00", -- $0e2b2
          58035 => x"00", -- $0e2b3
          58036 => x"00", -- $0e2b4
          58037 => x"00", -- $0e2b5
          58038 => x"00", -- $0e2b6
          58039 => x"00", -- $0e2b7
          58040 => x"00", -- $0e2b8
          58041 => x"00", -- $0e2b9
          58042 => x"00", -- $0e2ba
          58043 => x"00", -- $0e2bb
          58044 => x"00", -- $0e2bc
          58045 => x"00", -- $0e2bd
          58046 => x"00", -- $0e2be
          58047 => x"00", -- $0e2bf
          58048 => x"00", -- $0e2c0
          58049 => x"00", -- $0e2c1
          58050 => x"00", -- $0e2c2
          58051 => x"00", -- $0e2c3
          58052 => x"00", -- $0e2c4
          58053 => x"00", -- $0e2c5
          58054 => x"00", -- $0e2c6
          58055 => x"00", -- $0e2c7
          58056 => x"00", -- $0e2c8
          58057 => x"00", -- $0e2c9
          58058 => x"00", -- $0e2ca
          58059 => x"00", -- $0e2cb
          58060 => x"00", -- $0e2cc
          58061 => x"00", -- $0e2cd
          58062 => x"00", -- $0e2ce
          58063 => x"00", -- $0e2cf
          58064 => x"00", -- $0e2d0
          58065 => x"00", -- $0e2d1
          58066 => x"00", -- $0e2d2
          58067 => x"00", -- $0e2d3
          58068 => x"00", -- $0e2d4
          58069 => x"00", -- $0e2d5
          58070 => x"00", -- $0e2d6
          58071 => x"00", -- $0e2d7
          58072 => x"00", -- $0e2d8
          58073 => x"00", -- $0e2d9
          58074 => x"00", -- $0e2da
          58075 => x"00", -- $0e2db
          58076 => x"00", -- $0e2dc
          58077 => x"00", -- $0e2dd
          58078 => x"00", -- $0e2de
          58079 => x"00", -- $0e2df
          58080 => x"00", -- $0e2e0
          58081 => x"00", -- $0e2e1
          58082 => x"00", -- $0e2e2
          58083 => x"00", -- $0e2e3
          58084 => x"00", -- $0e2e4
          58085 => x"00", -- $0e2e5
          58086 => x"00", -- $0e2e6
          58087 => x"00", -- $0e2e7
          58088 => x"00", -- $0e2e8
          58089 => x"00", -- $0e2e9
          58090 => x"00", -- $0e2ea
          58091 => x"00", -- $0e2eb
          58092 => x"00", -- $0e2ec
          58093 => x"00", -- $0e2ed
          58094 => x"00", -- $0e2ee
          58095 => x"00", -- $0e2ef
          58096 => x"00", -- $0e2f0
          58097 => x"00", -- $0e2f1
          58098 => x"00", -- $0e2f2
          58099 => x"00", -- $0e2f3
          58100 => x"00", -- $0e2f4
          58101 => x"00", -- $0e2f5
          58102 => x"00", -- $0e2f6
          58103 => x"00", -- $0e2f7
          58104 => x"00", -- $0e2f8
          58105 => x"00", -- $0e2f9
          58106 => x"00", -- $0e2fa
          58107 => x"00", -- $0e2fb
          58108 => x"00", -- $0e2fc
          58109 => x"00", -- $0e2fd
          58110 => x"00", -- $0e2fe
          58111 => x"00", -- $0e2ff
          58112 => x"00", -- $0e300
          58113 => x"00", -- $0e301
          58114 => x"00", -- $0e302
          58115 => x"00", -- $0e303
          58116 => x"00", -- $0e304
          58117 => x"00", -- $0e305
          58118 => x"00", -- $0e306
          58119 => x"00", -- $0e307
          58120 => x"00", -- $0e308
          58121 => x"00", -- $0e309
          58122 => x"00", -- $0e30a
          58123 => x"00", -- $0e30b
          58124 => x"00", -- $0e30c
          58125 => x"00", -- $0e30d
          58126 => x"00", -- $0e30e
          58127 => x"00", -- $0e30f
          58128 => x"00", -- $0e310
          58129 => x"00", -- $0e311
          58130 => x"00", -- $0e312
          58131 => x"00", -- $0e313
          58132 => x"00", -- $0e314
          58133 => x"00", -- $0e315
          58134 => x"00", -- $0e316
          58135 => x"00", -- $0e317
          58136 => x"00", -- $0e318
          58137 => x"00", -- $0e319
          58138 => x"00", -- $0e31a
          58139 => x"00", -- $0e31b
          58140 => x"00", -- $0e31c
          58141 => x"00", -- $0e31d
          58142 => x"00", -- $0e31e
          58143 => x"00", -- $0e31f
          58144 => x"00", -- $0e320
          58145 => x"00", -- $0e321
          58146 => x"00", -- $0e322
          58147 => x"00", -- $0e323
          58148 => x"00", -- $0e324
          58149 => x"00", -- $0e325
          58150 => x"00", -- $0e326
          58151 => x"00", -- $0e327
          58152 => x"00", -- $0e328
          58153 => x"00", -- $0e329
          58154 => x"00", -- $0e32a
          58155 => x"00", -- $0e32b
          58156 => x"00", -- $0e32c
          58157 => x"00", -- $0e32d
          58158 => x"00", -- $0e32e
          58159 => x"00", -- $0e32f
          58160 => x"00", -- $0e330
          58161 => x"00", -- $0e331
          58162 => x"00", -- $0e332
          58163 => x"00", -- $0e333
          58164 => x"00", -- $0e334
          58165 => x"00", -- $0e335
          58166 => x"00", -- $0e336
          58167 => x"00", -- $0e337
          58168 => x"00", -- $0e338
          58169 => x"00", -- $0e339
          58170 => x"00", -- $0e33a
          58171 => x"00", -- $0e33b
          58172 => x"00", -- $0e33c
          58173 => x"00", -- $0e33d
          58174 => x"00", -- $0e33e
          58175 => x"00", -- $0e33f
          58176 => x"00", -- $0e340
          58177 => x"00", -- $0e341
          58178 => x"00", -- $0e342
          58179 => x"00", -- $0e343
          58180 => x"00", -- $0e344
          58181 => x"00", -- $0e345
          58182 => x"00", -- $0e346
          58183 => x"00", -- $0e347
          58184 => x"00", -- $0e348
          58185 => x"00", -- $0e349
          58186 => x"00", -- $0e34a
          58187 => x"00", -- $0e34b
          58188 => x"00", -- $0e34c
          58189 => x"00", -- $0e34d
          58190 => x"00", -- $0e34e
          58191 => x"00", -- $0e34f
          58192 => x"00", -- $0e350
          58193 => x"00", -- $0e351
          58194 => x"00", -- $0e352
          58195 => x"00", -- $0e353
          58196 => x"00", -- $0e354
          58197 => x"00", -- $0e355
          58198 => x"00", -- $0e356
          58199 => x"00", -- $0e357
          58200 => x"00", -- $0e358
          58201 => x"00", -- $0e359
          58202 => x"00", -- $0e35a
          58203 => x"00", -- $0e35b
          58204 => x"00", -- $0e35c
          58205 => x"00", -- $0e35d
          58206 => x"00", -- $0e35e
          58207 => x"00", -- $0e35f
          58208 => x"00", -- $0e360
          58209 => x"00", -- $0e361
          58210 => x"00", -- $0e362
          58211 => x"00", -- $0e363
          58212 => x"00", -- $0e364
          58213 => x"00", -- $0e365
          58214 => x"00", -- $0e366
          58215 => x"00", -- $0e367
          58216 => x"00", -- $0e368
          58217 => x"00", -- $0e369
          58218 => x"00", -- $0e36a
          58219 => x"00", -- $0e36b
          58220 => x"00", -- $0e36c
          58221 => x"00", -- $0e36d
          58222 => x"00", -- $0e36e
          58223 => x"00", -- $0e36f
          58224 => x"00", -- $0e370
          58225 => x"00", -- $0e371
          58226 => x"00", -- $0e372
          58227 => x"00", -- $0e373
          58228 => x"00", -- $0e374
          58229 => x"00", -- $0e375
          58230 => x"00", -- $0e376
          58231 => x"00", -- $0e377
          58232 => x"00", -- $0e378
          58233 => x"00", -- $0e379
          58234 => x"00", -- $0e37a
          58235 => x"00", -- $0e37b
          58236 => x"00", -- $0e37c
          58237 => x"00", -- $0e37d
          58238 => x"00", -- $0e37e
          58239 => x"00", -- $0e37f
          58240 => x"00", -- $0e380
          58241 => x"00", -- $0e381
          58242 => x"00", -- $0e382
          58243 => x"00", -- $0e383
          58244 => x"00", -- $0e384
          58245 => x"00", -- $0e385
          58246 => x"00", -- $0e386
          58247 => x"00", -- $0e387
          58248 => x"00", -- $0e388
          58249 => x"00", -- $0e389
          58250 => x"00", -- $0e38a
          58251 => x"00", -- $0e38b
          58252 => x"00", -- $0e38c
          58253 => x"00", -- $0e38d
          58254 => x"00", -- $0e38e
          58255 => x"00", -- $0e38f
          58256 => x"00", -- $0e390
          58257 => x"00", -- $0e391
          58258 => x"00", -- $0e392
          58259 => x"00", -- $0e393
          58260 => x"00", -- $0e394
          58261 => x"00", -- $0e395
          58262 => x"00", -- $0e396
          58263 => x"00", -- $0e397
          58264 => x"00", -- $0e398
          58265 => x"00", -- $0e399
          58266 => x"00", -- $0e39a
          58267 => x"00", -- $0e39b
          58268 => x"00", -- $0e39c
          58269 => x"00", -- $0e39d
          58270 => x"00", -- $0e39e
          58271 => x"00", -- $0e39f
          58272 => x"00", -- $0e3a0
          58273 => x"00", -- $0e3a1
          58274 => x"00", -- $0e3a2
          58275 => x"00", -- $0e3a3
          58276 => x"00", -- $0e3a4
          58277 => x"00", -- $0e3a5
          58278 => x"00", -- $0e3a6
          58279 => x"00", -- $0e3a7
          58280 => x"00", -- $0e3a8
          58281 => x"00", -- $0e3a9
          58282 => x"00", -- $0e3aa
          58283 => x"00", -- $0e3ab
          58284 => x"00", -- $0e3ac
          58285 => x"00", -- $0e3ad
          58286 => x"00", -- $0e3ae
          58287 => x"00", -- $0e3af
          58288 => x"00", -- $0e3b0
          58289 => x"00", -- $0e3b1
          58290 => x"00", -- $0e3b2
          58291 => x"00", -- $0e3b3
          58292 => x"00", -- $0e3b4
          58293 => x"00", -- $0e3b5
          58294 => x"00", -- $0e3b6
          58295 => x"00", -- $0e3b7
          58296 => x"00", -- $0e3b8
          58297 => x"00", -- $0e3b9
          58298 => x"00", -- $0e3ba
          58299 => x"00", -- $0e3bb
          58300 => x"00", -- $0e3bc
          58301 => x"00", -- $0e3bd
          58302 => x"00", -- $0e3be
          58303 => x"00", -- $0e3bf
          58304 => x"00", -- $0e3c0
          58305 => x"00", -- $0e3c1
          58306 => x"00", -- $0e3c2
          58307 => x"00", -- $0e3c3
          58308 => x"00", -- $0e3c4
          58309 => x"00", -- $0e3c5
          58310 => x"00", -- $0e3c6
          58311 => x"00", -- $0e3c7
          58312 => x"00", -- $0e3c8
          58313 => x"00", -- $0e3c9
          58314 => x"00", -- $0e3ca
          58315 => x"00", -- $0e3cb
          58316 => x"00", -- $0e3cc
          58317 => x"00", -- $0e3cd
          58318 => x"00", -- $0e3ce
          58319 => x"00", -- $0e3cf
          58320 => x"00", -- $0e3d0
          58321 => x"00", -- $0e3d1
          58322 => x"00", -- $0e3d2
          58323 => x"00", -- $0e3d3
          58324 => x"00", -- $0e3d4
          58325 => x"00", -- $0e3d5
          58326 => x"00", -- $0e3d6
          58327 => x"00", -- $0e3d7
          58328 => x"00", -- $0e3d8
          58329 => x"00", -- $0e3d9
          58330 => x"00", -- $0e3da
          58331 => x"00", -- $0e3db
          58332 => x"00", -- $0e3dc
          58333 => x"00", -- $0e3dd
          58334 => x"00", -- $0e3de
          58335 => x"00", -- $0e3df
          58336 => x"00", -- $0e3e0
          58337 => x"00", -- $0e3e1
          58338 => x"00", -- $0e3e2
          58339 => x"00", -- $0e3e3
          58340 => x"00", -- $0e3e4
          58341 => x"00", -- $0e3e5
          58342 => x"00", -- $0e3e6
          58343 => x"00", -- $0e3e7
          58344 => x"00", -- $0e3e8
          58345 => x"00", -- $0e3e9
          58346 => x"00", -- $0e3ea
          58347 => x"00", -- $0e3eb
          58348 => x"00", -- $0e3ec
          58349 => x"00", -- $0e3ed
          58350 => x"00", -- $0e3ee
          58351 => x"00", -- $0e3ef
          58352 => x"00", -- $0e3f0
          58353 => x"00", -- $0e3f1
          58354 => x"00", -- $0e3f2
          58355 => x"00", -- $0e3f3
          58356 => x"00", -- $0e3f4
          58357 => x"00", -- $0e3f5
          58358 => x"00", -- $0e3f6
          58359 => x"00", -- $0e3f7
          58360 => x"00", -- $0e3f8
          58361 => x"00", -- $0e3f9
          58362 => x"00", -- $0e3fa
          58363 => x"00", -- $0e3fb
          58364 => x"00", -- $0e3fc
          58365 => x"00", -- $0e3fd
          58366 => x"00", -- $0e3fe
          58367 => x"00", -- $0e3ff
          58368 => x"00", -- $0e400
          58369 => x"00", -- $0e401
          58370 => x"00", -- $0e402
          58371 => x"00", -- $0e403
          58372 => x"00", -- $0e404
          58373 => x"00", -- $0e405
          58374 => x"00", -- $0e406
          58375 => x"00", -- $0e407
          58376 => x"00", -- $0e408
          58377 => x"00", -- $0e409
          58378 => x"00", -- $0e40a
          58379 => x"00", -- $0e40b
          58380 => x"00", -- $0e40c
          58381 => x"00", -- $0e40d
          58382 => x"00", -- $0e40e
          58383 => x"00", -- $0e40f
          58384 => x"00", -- $0e410
          58385 => x"00", -- $0e411
          58386 => x"00", -- $0e412
          58387 => x"00", -- $0e413
          58388 => x"00", -- $0e414
          58389 => x"00", -- $0e415
          58390 => x"00", -- $0e416
          58391 => x"00", -- $0e417
          58392 => x"00", -- $0e418
          58393 => x"00", -- $0e419
          58394 => x"00", -- $0e41a
          58395 => x"00", -- $0e41b
          58396 => x"00", -- $0e41c
          58397 => x"00", -- $0e41d
          58398 => x"00", -- $0e41e
          58399 => x"00", -- $0e41f
          58400 => x"00", -- $0e420
          58401 => x"00", -- $0e421
          58402 => x"00", -- $0e422
          58403 => x"00", -- $0e423
          58404 => x"00", -- $0e424
          58405 => x"00", -- $0e425
          58406 => x"00", -- $0e426
          58407 => x"00", -- $0e427
          58408 => x"00", -- $0e428
          58409 => x"00", -- $0e429
          58410 => x"00", -- $0e42a
          58411 => x"00", -- $0e42b
          58412 => x"00", -- $0e42c
          58413 => x"00", -- $0e42d
          58414 => x"00", -- $0e42e
          58415 => x"00", -- $0e42f
          58416 => x"00", -- $0e430
          58417 => x"00", -- $0e431
          58418 => x"00", -- $0e432
          58419 => x"00", -- $0e433
          58420 => x"00", -- $0e434
          58421 => x"00", -- $0e435
          58422 => x"00", -- $0e436
          58423 => x"00", -- $0e437
          58424 => x"00", -- $0e438
          58425 => x"00", -- $0e439
          58426 => x"00", -- $0e43a
          58427 => x"00", -- $0e43b
          58428 => x"00", -- $0e43c
          58429 => x"00", -- $0e43d
          58430 => x"00", -- $0e43e
          58431 => x"00", -- $0e43f
          58432 => x"00", -- $0e440
          58433 => x"00", -- $0e441
          58434 => x"00", -- $0e442
          58435 => x"00", -- $0e443
          58436 => x"00", -- $0e444
          58437 => x"00", -- $0e445
          58438 => x"00", -- $0e446
          58439 => x"00", -- $0e447
          58440 => x"00", -- $0e448
          58441 => x"00", -- $0e449
          58442 => x"00", -- $0e44a
          58443 => x"00", -- $0e44b
          58444 => x"00", -- $0e44c
          58445 => x"00", -- $0e44d
          58446 => x"00", -- $0e44e
          58447 => x"00", -- $0e44f
          58448 => x"00", -- $0e450
          58449 => x"00", -- $0e451
          58450 => x"00", -- $0e452
          58451 => x"00", -- $0e453
          58452 => x"00", -- $0e454
          58453 => x"00", -- $0e455
          58454 => x"00", -- $0e456
          58455 => x"00", -- $0e457
          58456 => x"00", -- $0e458
          58457 => x"00", -- $0e459
          58458 => x"00", -- $0e45a
          58459 => x"00", -- $0e45b
          58460 => x"00", -- $0e45c
          58461 => x"00", -- $0e45d
          58462 => x"00", -- $0e45e
          58463 => x"00", -- $0e45f
          58464 => x"00", -- $0e460
          58465 => x"00", -- $0e461
          58466 => x"00", -- $0e462
          58467 => x"00", -- $0e463
          58468 => x"00", -- $0e464
          58469 => x"00", -- $0e465
          58470 => x"00", -- $0e466
          58471 => x"00", -- $0e467
          58472 => x"00", -- $0e468
          58473 => x"00", -- $0e469
          58474 => x"00", -- $0e46a
          58475 => x"00", -- $0e46b
          58476 => x"00", -- $0e46c
          58477 => x"00", -- $0e46d
          58478 => x"00", -- $0e46e
          58479 => x"00", -- $0e46f
          58480 => x"00", -- $0e470
          58481 => x"00", -- $0e471
          58482 => x"00", -- $0e472
          58483 => x"00", -- $0e473
          58484 => x"00", -- $0e474
          58485 => x"00", -- $0e475
          58486 => x"00", -- $0e476
          58487 => x"00", -- $0e477
          58488 => x"00", -- $0e478
          58489 => x"00", -- $0e479
          58490 => x"00", -- $0e47a
          58491 => x"00", -- $0e47b
          58492 => x"00", -- $0e47c
          58493 => x"00", -- $0e47d
          58494 => x"00", -- $0e47e
          58495 => x"00", -- $0e47f
          58496 => x"00", -- $0e480
          58497 => x"00", -- $0e481
          58498 => x"00", -- $0e482
          58499 => x"00", -- $0e483
          58500 => x"00", -- $0e484
          58501 => x"00", -- $0e485
          58502 => x"00", -- $0e486
          58503 => x"00", -- $0e487
          58504 => x"00", -- $0e488
          58505 => x"00", -- $0e489
          58506 => x"00", -- $0e48a
          58507 => x"00", -- $0e48b
          58508 => x"00", -- $0e48c
          58509 => x"00", -- $0e48d
          58510 => x"00", -- $0e48e
          58511 => x"00", -- $0e48f
          58512 => x"00", -- $0e490
          58513 => x"00", -- $0e491
          58514 => x"00", -- $0e492
          58515 => x"00", -- $0e493
          58516 => x"00", -- $0e494
          58517 => x"00", -- $0e495
          58518 => x"00", -- $0e496
          58519 => x"00", -- $0e497
          58520 => x"00", -- $0e498
          58521 => x"00", -- $0e499
          58522 => x"00", -- $0e49a
          58523 => x"00", -- $0e49b
          58524 => x"00", -- $0e49c
          58525 => x"00", -- $0e49d
          58526 => x"00", -- $0e49e
          58527 => x"00", -- $0e49f
          58528 => x"00", -- $0e4a0
          58529 => x"00", -- $0e4a1
          58530 => x"00", -- $0e4a2
          58531 => x"00", -- $0e4a3
          58532 => x"00", -- $0e4a4
          58533 => x"00", -- $0e4a5
          58534 => x"00", -- $0e4a6
          58535 => x"00", -- $0e4a7
          58536 => x"00", -- $0e4a8
          58537 => x"00", -- $0e4a9
          58538 => x"00", -- $0e4aa
          58539 => x"00", -- $0e4ab
          58540 => x"00", -- $0e4ac
          58541 => x"00", -- $0e4ad
          58542 => x"00", -- $0e4ae
          58543 => x"00", -- $0e4af
          58544 => x"00", -- $0e4b0
          58545 => x"00", -- $0e4b1
          58546 => x"00", -- $0e4b2
          58547 => x"00", -- $0e4b3
          58548 => x"00", -- $0e4b4
          58549 => x"00", -- $0e4b5
          58550 => x"00", -- $0e4b6
          58551 => x"00", -- $0e4b7
          58552 => x"00", -- $0e4b8
          58553 => x"00", -- $0e4b9
          58554 => x"00", -- $0e4ba
          58555 => x"00", -- $0e4bb
          58556 => x"00", -- $0e4bc
          58557 => x"00", -- $0e4bd
          58558 => x"00", -- $0e4be
          58559 => x"00", -- $0e4bf
          58560 => x"00", -- $0e4c0
          58561 => x"00", -- $0e4c1
          58562 => x"00", -- $0e4c2
          58563 => x"00", -- $0e4c3
          58564 => x"00", -- $0e4c4
          58565 => x"00", -- $0e4c5
          58566 => x"00", -- $0e4c6
          58567 => x"00", -- $0e4c7
          58568 => x"00", -- $0e4c8
          58569 => x"00", -- $0e4c9
          58570 => x"00", -- $0e4ca
          58571 => x"00", -- $0e4cb
          58572 => x"00", -- $0e4cc
          58573 => x"00", -- $0e4cd
          58574 => x"00", -- $0e4ce
          58575 => x"00", -- $0e4cf
          58576 => x"00", -- $0e4d0
          58577 => x"00", -- $0e4d1
          58578 => x"00", -- $0e4d2
          58579 => x"00", -- $0e4d3
          58580 => x"00", -- $0e4d4
          58581 => x"00", -- $0e4d5
          58582 => x"00", -- $0e4d6
          58583 => x"00", -- $0e4d7
          58584 => x"00", -- $0e4d8
          58585 => x"00", -- $0e4d9
          58586 => x"00", -- $0e4da
          58587 => x"00", -- $0e4db
          58588 => x"00", -- $0e4dc
          58589 => x"00", -- $0e4dd
          58590 => x"00", -- $0e4de
          58591 => x"00", -- $0e4df
          58592 => x"00", -- $0e4e0
          58593 => x"00", -- $0e4e1
          58594 => x"00", -- $0e4e2
          58595 => x"00", -- $0e4e3
          58596 => x"00", -- $0e4e4
          58597 => x"00", -- $0e4e5
          58598 => x"00", -- $0e4e6
          58599 => x"00", -- $0e4e7
          58600 => x"00", -- $0e4e8
          58601 => x"00", -- $0e4e9
          58602 => x"00", -- $0e4ea
          58603 => x"00", -- $0e4eb
          58604 => x"00", -- $0e4ec
          58605 => x"00", -- $0e4ed
          58606 => x"00", -- $0e4ee
          58607 => x"00", -- $0e4ef
          58608 => x"00", -- $0e4f0
          58609 => x"00", -- $0e4f1
          58610 => x"00", -- $0e4f2
          58611 => x"00", -- $0e4f3
          58612 => x"00", -- $0e4f4
          58613 => x"00", -- $0e4f5
          58614 => x"00", -- $0e4f6
          58615 => x"00", -- $0e4f7
          58616 => x"00", -- $0e4f8
          58617 => x"00", -- $0e4f9
          58618 => x"00", -- $0e4fa
          58619 => x"00", -- $0e4fb
          58620 => x"00", -- $0e4fc
          58621 => x"00", -- $0e4fd
          58622 => x"00", -- $0e4fe
          58623 => x"00", -- $0e4ff
          58624 => x"00", -- $0e500
          58625 => x"00", -- $0e501
          58626 => x"00", -- $0e502
          58627 => x"00", -- $0e503
          58628 => x"00", -- $0e504
          58629 => x"00", -- $0e505
          58630 => x"00", -- $0e506
          58631 => x"00", -- $0e507
          58632 => x"00", -- $0e508
          58633 => x"00", -- $0e509
          58634 => x"00", -- $0e50a
          58635 => x"00", -- $0e50b
          58636 => x"00", -- $0e50c
          58637 => x"00", -- $0e50d
          58638 => x"00", -- $0e50e
          58639 => x"00", -- $0e50f
          58640 => x"00", -- $0e510
          58641 => x"00", -- $0e511
          58642 => x"00", -- $0e512
          58643 => x"00", -- $0e513
          58644 => x"00", -- $0e514
          58645 => x"00", -- $0e515
          58646 => x"00", -- $0e516
          58647 => x"00", -- $0e517
          58648 => x"00", -- $0e518
          58649 => x"00", -- $0e519
          58650 => x"00", -- $0e51a
          58651 => x"00", -- $0e51b
          58652 => x"00", -- $0e51c
          58653 => x"00", -- $0e51d
          58654 => x"00", -- $0e51e
          58655 => x"00", -- $0e51f
          58656 => x"00", -- $0e520
          58657 => x"00", -- $0e521
          58658 => x"00", -- $0e522
          58659 => x"00", -- $0e523
          58660 => x"00", -- $0e524
          58661 => x"00", -- $0e525
          58662 => x"00", -- $0e526
          58663 => x"00", -- $0e527
          58664 => x"00", -- $0e528
          58665 => x"00", -- $0e529
          58666 => x"00", -- $0e52a
          58667 => x"00", -- $0e52b
          58668 => x"00", -- $0e52c
          58669 => x"00", -- $0e52d
          58670 => x"00", -- $0e52e
          58671 => x"00", -- $0e52f
          58672 => x"00", -- $0e530
          58673 => x"00", -- $0e531
          58674 => x"00", -- $0e532
          58675 => x"00", -- $0e533
          58676 => x"00", -- $0e534
          58677 => x"00", -- $0e535
          58678 => x"00", -- $0e536
          58679 => x"00", -- $0e537
          58680 => x"00", -- $0e538
          58681 => x"00", -- $0e539
          58682 => x"00", -- $0e53a
          58683 => x"00", -- $0e53b
          58684 => x"00", -- $0e53c
          58685 => x"00", -- $0e53d
          58686 => x"00", -- $0e53e
          58687 => x"00", -- $0e53f
          58688 => x"00", -- $0e540
          58689 => x"00", -- $0e541
          58690 => x"00", -- $0e542
          58691 => x"00", -- $0e543
          58692 => x"00", -- $0e544
          58693 => x"00", -- $0e545
          58694 => x"00", -- $0e546
          58695 => x"00", -- $0e547
          58696 => x"00", -- $0e548
          58697 => x"00", -- $0e549
          58698 => x"00", -- $0e54a
          58699 => x"00", -- $0e54b
          58700 => x"00", -- $0e54c
          58701 => x"00", -- $0e54d
          58702 => x"00", -- $0e54e
          58703 => x"00", -- $0e54f
          58704 => x"00", -- $0e550
          58705 => x"00", -- $0e551
          58706 => x"00", -- $0e552
          58707 => x"00", -- $0e553
          58708 => x"00", -- $0e554
          58709 => x"00", -- $0e555
          58710 => x"00", -- $0e556
          58711 => x"00", -- $0e557
          58712 => x"00", -- $0e558
          58713 => x"00", -- $0e559
          58714 => x"00", -- $0e55a
          58715 => x"00", -- $0e55b
          58716 => x"00", -- $0e55c
          58717 => x"00", -- $0e55d
          58718 => x"00", -- $0e55e
          58719 => x"00", -- $0e55f
          58720 => x"00", -- $0e560
          58721 => x"00", -- $0e561
          58722 => x"00", -- $0e562
          58723 => x"00", -- $0e563
          58724 => x"00", -- $0e564
          58725 => x"00", -- $0e565
          58726 => x"00", -- $0e566
          58727 => x"00", -- $0e567
          58728 => x"00", -- $0e568
          58729 => x"00", -- $0e569
          58730 => x"00", -- $0e56a
          58731 => x"00", -- $0e56b
          58732 => x"00", -- $0e56c
          58733 => x"00", -- $0e56d
          58734 => x"00", -- $0e56e
          58735 => x"00", -- $0e56f
          58736 => x"00", -- $0e570
          58737 => x"00", -- $0e571
          58738 => x"00", -- $0e572
          58739 => x"00", -- $0e573
          58740 => x"00", -- $0e574
          58741 => x"00", -- $0e575
          58742 => x"00", -- $0e576
          58743 => x"00", -- $0e577
          58744 => x"00", -- $0e578
          58745 => x"00", -- $0e579
          58746 => x"00", -- $0e57a
          58747 => x"00", -- $0e57b
          58748 => x"00", -- $0e57c
          58749 => x"00", -- $0e57d
          58750 => x"00", -- $0e57e
          58751 => x"00", -- $0e57f
          58752 => x"00", -- $0e580
          58753 => x"00", -- $0e581
          58754 => x"00", -- $0e582
          58755 => x"00", -- $0e583
          58756 => x"00", -- $0e584
          58757 => x"00", -- $0e585
          58758 => x"00", -- $0e586
          58759 => x"00", -- $0e587
          58760 => x"00", -- $0e588
          58761 => x"00", -- $0e589
          58762 => x"00", -- $0e58a
          58763 => x"00", -- $0e58b
          58764 => x"00", -- $0e58c
          58765 => x"00", -- $0e58d
          58766 => x"00", -- $0e58e
          58767 => x"00", -- $0e58f
          58768 => x"00", -- $0e590
          58769 => x"00", -- $0e591
          58770 => x"00", -- $0e592
          58771 => x"00", -- $0e593
          58772 => x"00", -- $0e594
          58773 => x"00", -- $0e595
          58774 => x"00", -- $0e596
          58775 => x"00", -- $0e597
          58776 => x"00", -- $0e598
          58777 => x"00", -- $0e599
          58778 => x"00", -- $0e59a
          58779 => x"00", -- $0e59b
          58780 => x"00", -- $0e59c
          58781 => x"00", -- $0e59d
          58782 => x"00", -- $0e59e
          58783 => x"00", -- $0e59f
          58784 => x"00", -- $0e5a0
          58785 => x"00", -- $0e5a1
          58786 => x"00", -- $0e5a2
          58787 => x"00", -- $0e5a3
          58788 => x"00", -- $0e5a4
          58789 => x"00", -- $0e5a5
          58790 => x"00", -- $0e5a6
          58791 => x"00", -- $0e5a7
          58792 => x"00", -- $0e5a8
          58793 => x"00", -- $0e5a9
          58794 => x"00", -- $0e5aa
          58795 => x"00", -- $0e5ab
          58796 => x"00", -- $0e5ac
          58797 => x"00", -- $0e5ad
          58798 => x"00", -- $0e5ae
          58799 => x"00", -- $0e5af
          58800 => x"00", -- $0e5b0
          58801 => x"00", -- $0e5b1
          58802 => x"00", -- $0e5b2
          58803 => x"00", -- $0e5b3
          58804 => x"00", -- $0e5b4
          58805 => x"00", -- $0e5b5
          58806 => x"00", -- $0e5b6
          58807 => x"00", -- $0e5b7
          58808 => x"00", -- $0e5b8
          58809 => x"00", -- $0e5b9
          58810 => x"00", -- $0e5ba
          58811 => x"00", -- $0e5bb
          58812 => x"00", -- $0e5bc
          58813 => x"00", -- $0e5bd
          58814 => x"00", -- $0e5be
          58815 => x"00", -- $0e5bf
          58816 => x"00", -- $0e5c0
          58817 => x"00", -- $0e5c1
          58818 => x"00", -- $0e5c2
          58819 => x"00", -- $0e5c3
          58820 => x"00", -- $0e5c4
          58821 => x"00", -- $0e5c5
          58822 => x"00", -- $0e5c6
          58823 => x"00", -- $0e5c7
          58824 => x"00", -- $0e5c8
          58825 => x"00", -- $0e5c9
          58826 => x"00", -- $0e5ca
          58827 => x"00", -- $0e5cb
          58828 => x"00", -- $0e5cc
          58829 => x"00", -- $0e5cd
          58830 => x"00", -- $0e5ce
          58831 => x"00", -- $0e5cf
          58832 => x"00", -- $0e5d0
          58833 => x"00", -- $0e5d1
          58834 => x"00", -- $0e5d2
          58835 => x"00", -- $0e5d3
          58836 => x"00", -- $0e5d4
          58837 => x"00", -- $0e5d5
          58838 => x"00", -- $0e5d6
          58839 => x"00", -- $0e5d7
          58840 => x"00", -- $0e5d8
          58841 => x"00", -- $0e5d9
          58842 => x"00", -- $0e5da
          58843 => x"00", -- $0e5db
          58844 => x"00", -- $0e5dc
          58845 => x"00", -- $0e5dd
          58846 => x"00", -- $0e5de
          58847 => x"00", -- $0e5df
          58848 => x"00", -- $0e5e0
          58849 => x"00", -- $0e5e1
          58850 => x"00", -- $0e5e2
          58851 => x"00", -- $0e5e3
          58852 => x"00", -- $0e5e4
          58853 => x"00", -- $0e5e5
          58854 => x"00", -- $0e5e6
          58855 => x"00", -- $0e5e7
          58856 => x"00", -- $0e5e8
          58857 => x"00", -- $0e5e9
          58858 => x"00", -- $0e5ea
          58859 => x"00", -- $0e5eb
          58860 => x"00", -- $0e5ec
          58861 => x"00", -- $0e5ed
          58862 => x"00", -- $0e5ee
          58863 => x"00", -- $0e5ef
          58864 => x"00", -- $0e5f0
          58865 => x"00", -- $0e5f1
          58866 => x"00", -- $0e5f2
          58867 => x"00", -- $0e5f3
          58868 => x"00", -- $0e5f4
          58869 => x"00", -- $0e5f5
          58870 => x"00", -- $0e5f6
          58871 => x"00", -- $0e5f7
          58872 => x"00", -- $0e5f8
          58873 => x"00", -- $0e5f9
          58874 => x"00", -- $0e5fa
          58875 => x"00", -- $0e5fb
          58876 => x"00", -- $0e5fc
          58877 => x"00", -- $0e5fd
          58878 => x"00", -- $0e5fe
          58879 => x"00", -- $0e5ff
          58880 => x"00", -- $0e600
          58881 => x"00", -- $0e601
          58882 => x"00", -- $0e602
          58883 => x"00", -- $0e603
          58884 => x"00", -- $0e604
          58885 => x"00", -- $0e605
          58886 => x"00", -- $0e606
          58887 => x"00", -- $0e607
          58888 => x"00", -- $0e608
          58889 => x"00", -- $0e609
          58890 => x"00", -- $0e60a
          58891 => x"00", -- $0e60b
          58892 => x"00", -- $0e60c
          58893 => x"00", -- $0e60d
          58894 => x"00", -- $0e60e
          58895 => x"00", -- $0e60f
          58896 => x"00", -- $0e610
          58897 => x"00", -- $0e611
          58898 => x"00", -- $0e612
          58899 => x"00", -- $0e613
          58900 => x"00", -- $0e614
          58901 => x"00", -- $0e615
          58902 => x"00", -- $0e616
          58903 => x"00", -- $0e617
          58904 => x"00", -- $0e618
          58905 => x"00", -- $0e619
          58906 => x"00", -- $0e61a
          58907 => x"00", -- $0e61b
          58908 => x"00", -- $0e61c
          58909 => x"00", -- $0e61d
          58910 => x"00", -- $0e61e
          58911 => x"00", -- $0e61f
          58912 => x"00", -- $0e620
          58913 => x"00", -- $0e621
          58914 => x"00", -- $0e622
          58915 => x"00", -- $0e623
          58916 => x"00", -- $0e624
          58917 => x"00", -- $0e625
          58918 => x"00", -- $0e626
          58919 => x"00", -- $0e627
          58920 => x"00", -- $0e628
          58921 => x"00", -- $0e629
          58922 => x"00", -- $0e62a
          58923 => x"00", -- $0e62b
          58924 => x"00", -- $0e62c
          58925 => x"00", -- $0e62d
          58926 => x"00", -- $0e62e
          58927 => x"00", -- $0e62f
          58928 => x"00", -- $0e630
          58929 => x"00", -- $0e631
          58930 => x"00", -- $0e632
          58931 => x"00", -- $0e633
          58932 => x"00", -- $0e634
          58933 => x"00", -- $0e635
          58934 => x"00", -- $0e636
          58935 => x"00", -- $0e637
          58936 => x"00", -- $0e638
          58937 => x"00", -- $0e639
          58938 => x"00", -- $0e63a
          58939 => x"00", -- $0e63b
          58940 => x"00", -- $0e63c
          58941 => x"00", -- $0e63d
          58942 => x"00", -- $0e63e
          58943 => x"00", -- $0e63f
          58944 => x"00", -- $0e640
          58945 => x"00", -- $0e641
          58946 => x"00", -- $0e642
          58947 => x"00", -- $0e643
          58948 => x"00", -- $0e644
          58949 => x"00", -- $0e645
          58950 => x"00", -- $0e646
          58951 => x"00", -- $0e647
          58952 => x"00", -- $0e648
          58953 => x"00", -- $0e649
          58954 => x"00", -- $0e64a
          58955 => x"00", -- $0e64b
          58956 => x"00", -- $0e64c
          58957 => x"00", -- $0e64d
          58958 => x"00", -- $0e64e
          58959 => x"00", -- $0e64f
          58960 => x"00", -- $0e650
          58961 => x"00", -- $0e651
          58962 => x"00", -- $0e652
          58963 => x"00", -- $0e653
          58964 => x"00", -- $0e654
          58965 => x"00", -- $0e655
          58966 => x"00", -- $0e656
          58967 => x"00", -- $0e657
          58968 => x"00", -- $0e658
          58969 => x"00", -- $0e659
          58970 => x"00", -- $0e65a
          58971 => x"00", -- $0e65b
          58972 => x"00", -- $0e65c
          58973 => x"00", -- $0e65d
          58974 => x"00", -- $0e65e
          58975 => x"00", -- $0e65f
          58976 => x"00", -- $0e660
          58977 => x"00", -- $0e661
          58978 => x"00", -- $0e662
          58979 => x"00", -- $0e663
          58980 => x"00", -- $0e664
          58981 => x"00", -- $0e665
          58982 => x"00", -- $0e666
          58983 => x"00", -- $0e667
          58984 => x"00", -- $0e668
          58985 => x"00", -- $0e669
          58986 => x"00", -- $0e66a
          58987 => x"00", -- $0e66b
          58988 => x"00", -- $0e66c
          58989 => x"00", -- $0e66d
          58990 => x"00", -- $0e66e
          58991 => x"00", -- $0e66f
          58992 => x"00", -- $0e670
          58993 => x"00", -- $0e671
          58994 => x"00", -- $0e672
          58995 => x"00", -- $0e673
          58996 => x"00", -- $0e674
          58997 => x"00", -- $0e675
          58998 => x"00", -- $0e676
          58999 => x"00", -- $0e677
          59000 => x"00", -- $0e678
          59001 => x"00", -- $0e679
          59002 => x"00", -- $0e67a
          59003 => x"00", -- $0e67b
          59004 => x"00", -- $0e67c
          59005 => x"00", -- $0e67d
          59006 => x"00", -- $0e67e
          59007 => x"00", -- $0e67f
          59008 => x"00", -- $0e680
          59009 => x"00", -- $0e681
          59010 => x"00", -- $0e682
          59011 => x"00", -- $0e683
          59012 => x"00", -- $0e684
          59013 => x"00", -- $0e685
          59014 => x"00", -- $0e686
          59015 => x"00", -- $0e687
          59016 => x"00", -- $0e688
          59017 => x"00", -- $0e689
          59018 => x"00", -- $0e68a
          59019 => x"00", -- $0e68b
          59020 => x"00", -- $0e68c
          59021 => x"00", -- $0e68d
          59022 => x"00", -- $0e68e
          59023 => x"00", -- $0e68f
          59024 => x"00", -- $0e690
          59025 => x"00", -- $0e691
          59026 => x"00", -- $0e692
          59027 => x"00", -- $0e693
          59028 => x"00", -- $0e694
          59029 => x"00", -- $0e695
          59030 => x"00", -- $0e696
          59031 => x"00", -- $0e697
          59032 => x"00", -- $0e698
          59033 => x"00", -- $0e699
          59034 => x"00", -- $0e69a
          59035 => x"00", -- $0e69b
          59036 => x"00", -- $0e69c
          59037 => x"00", -- $0e69d
          59038 => x"00", -- $0e69e
          59039 => x"00", -- $0e69f
          59040 => x"00", -- $0e6a0
          59041 => x"00", -- $0e6a1
          59042 => x"00", -- $0e6a2
          59043 => x"00", -- $0e6a3
          59044 => x"00", -- $0e6a4
          59045 => x"00", -- $0e6a5
          59046 => x"00", -- $0e6a6
          59047 => x"00", -- $0e6a7
          59048 => x"00", -- $0e6a8
          59049 => x"00", -- $0e6a9
          59050 => x"00", -- $0e6aa
          59051 => x"00", -- $0e6ab
          59052 => x"00", -- $0e6ac
          59053 => x"00", -- $0e6ad
          59054 => x"00", -- $0e6ae
          59055 => x"00", -- $0e6af
          59056 => x"00", -- $0e6b0
          59057 => x"00", -- $0e6b1
          59058 => x"00", -- $0e6b2
          59059 => x"00", -- $0e6b3
          59060 => x"00", -- $0e6b4
          59061 => x"00", -- $0e6b5
          59062 => x"00", -- $0e6b6
          59063 => x"00", -- $0e6b7
          59064 => x"00", -- $0e6b8
          59065 => x"00", -- $0e6b9
          59066 => x"00", -- $0e6ba
          59067 => x"00", -- $0e6bb
          59068 => x"00", -- $0e6bc
          59069 => x"00", -- $0e6bd
          59070 => x"00", -- $0e6be
          59071 => x"00", -- $0e6bf
          59072 => x"00", -- $0e6c0
          59073 => x"00", -- $0e6c1
          59074 => x"00", -- $0e6c2
          59075 => x"00", -- $0e6c3
          59076 => x"00", -- $0e6c4
          59077 => x"00", -- $0e6c5
          59078 => x"00", -- $0e6c6
          59079 => x"00", -- $0e6c7
          59080 => x"00", -- $0e6c8
          59081 => x"00", -- $0e6c9
          59082 => x"00", -- $0e6ca
          59083 => x"00", -- $0e6cb
          59084 => x"00", -- $0e6cc
          59085 => x"00", -- $0e6cd
          59086 => x"00", -- $0e6ce
          59087 => x"00", -- $0e6cf
          59088 => x"00", -- $0e6d0
          59089 => x"00", -- $0e6d1
          59090 => x"00", -- $0e6d2
          59091 => x"00", -- $0e6d3
          59092 => x"00", -- $0e6d4
          59093 => x"00", -- $0e6d5
          59094 => x"00", -- $0e6d6
          59095 => x"00", -- $0e6d7
          59096 => x"00", -- $0e6d8
          59097 => x"00", -- $0e6d9
          59098 => x"00", -- $0e6da
          59099 => x"00", -- $0e6db
          59100 => x"00", -- $0e6dc
          59101 => x"00", -- $0e6dd
          59102 => x"00", -- $0e6de
          59103 => x"00", -- $0e6df
          59104 => x"00", -- $0e6e0
          59105 => x"00", -- $0e6e1
          59106 => x"00", -- $0e6e2
          59107 => x"00", -- $0e6e3
          59108 => x"00", -- $0e6e4
          59109 => x"00", -- $0e6e5
          59110 => x"00", -- $0e6e6
          59111 => x"00", -- $0e6e7
          59112 => x"00", -- $0e6e8
          59113 => x"00", -- $0e6e9
          59114 => x"00", -- $0e6ea
          59115 => x"00", -- $0e6eb
          59116 => x"00", -- $0e6ec
          59117 => x"00", -- $0e6ed
          59118 => x"00", -- $0e6ee
          59119 => x"00", -- $0e6ef
          59120 => x"00", -- $0e6f0
          59121 => x"00", -- $0e6f1
          59122 => x"00", -- $0e6f2
          59123 => x"00", -- $0e6f3
          59124 => x"00", -- $0e6f4
          59125 => x"00", -- $0e6f5
          59126 => x"00", -- $0e6f6
          59127 => x"00", -- $0e6f7
          59128 => x"00", -- $0e6f8
          59129 => x"00", -- $0e6f9
          59130 => x"00", -- $0e6fa
          59131 => x"00", -- $0e6fb
          59132 => x"00", -- $0e6fc
          59133 => x"00", -- $0e6fd
          59134 => x"00", -- $0e6fe
          59135 => x"00", -- $0e6ff
          59136 => x"00", -- $0e700
          59137 => x"00", -- $0e701
          59138 => x"00", -- $0e702
          59139 => x"00", -- $0e703
          59140 => x"00", -- $0e704
          59141 => x"00", -- $0e705
          59142 => x"00", -- $0e706
          59143 => x"00", -- $0e707
          59144 => x"00", -- $0e708
          59145 => x"00", -- $0e709
          59146 => x"00", -- $0e70a
          59147 => x"00", -- $0e70b
          59148 => x"00", -- $0e70c
          59149 => x"00", -- $0e70d
          59150 => x"00", -- $0e70e
          59151 => x"00", -- $0e70f
          59152 => x"00", -- $0e710
          59153 => x"00", -- $0e711
          59154 => x"00", -- $0e712
          59155 => x"00", -- $0e713
          59156 => x"00", -- $0e714
          59157 => x"00", -- $0e715
          59158 => x"00", -- $0e716
          59159 => x"00", -- $0e717
          59160 => x"00", -- $0e718
          59161 => x"00", -- $0e719
          59162 => x"00", -- $0e71a
          59163 => x"00", -- $0e71b
          59164 => x"00", -- $0e71c
          59165 => x"00", -- $0e71d
          59166 => x"00", -- $0e71e
          59167 => x"00", -- $0e71f
          59168 => x"00", -- $0e720
          59169 => x"00", -- $0e721
          59170 => x"00", -- $0e722
          59171 => x"00", -- $0e723
          59172 => x"00", -- $0e724
          59173 => x"00", -- $0e725
          59174 => x"00", -- $0e726
          59175 => x"00", -- $0e727
          59176 => x"00", -- $0e728
          59177 => x"00", -- $0e729
          59178 => x"00", -- $0e72a
          59179 => x"00", -- $0e72b
          59180 => x"00", -- $0e72c
          59181 => x"00", -- $0e72d
          59182 => x"00", -- $0e72e
          59183 => x"00", -- $0e72f
          59184 => x"00", -- $0e730
          59185 => x"00", -- $0e731
          59186 => x"00", -- $0e732
          59187 => x"00", -- $0e733
          59188 => x"00", -- $0e734
          59189 => x"00", -- $0e735
          59190 => x"00", -- $0e736
          59191 => x"00", -- $0e737
          59192 => x"00", -- $0e738
          59193 => x"00", -- $0e739
          59194 => x"00", -- $0e73a
          59195 => x"00", -- $0e73b
          59196 => x"00", -- $0e73c
          59197 => x"00", -- $0e73d
          59198 => x"00", -- $0e73e
          59199 => x"00", -- $0e73f
          59200 => x"00", -- $0e740
          59201 => x"00", -- $0e741
          59202 => x"00", -- $0e742
          59203 => x"00", -- $0e743
          59204 => x"00", -- $0e744
          59205 => x"00", -- $0e745
          59206 => x"00", -- $0e746
          59207 => x"00", -- $0e747
          59208 => x"00", -- $0e748
          59209 => x"00", -- $0e749
          59210 => x"00", -- $0e74a
          59211 => x"00", -- $0e74b
          59212 => x"00", -- $0e74c
          59213 => x"00", -- $0e74d
          59214 => x"00", -- $0e74e
          59215 => x"00", -- $0e74f
          59216 => x"00", -- $0e750
          59217 => x"00", -- $0e751
          59218 => x"00", -- $0e752
          59219 => x"00", -- $0e753
          59220 => x"00", -- $0e754
          59221 => x"00", -- $0e755
          59222 => x"00", -- $0e756
          59223 => x"00", -- $0e757
          59224 => x"00", -- $0e758
          59225 => x"00", -- $0e759
          59226 => x"00", -- $0e75a
          59227 => x"00", -- $0e75b
          59228 => x"00", -- $0e75c
          59229 => x"00", -- $0e75d
          59230 => x"00", -- $0e75e
          59231 => x"00", -- $0e75f
          59232 => x"00", -- $0e760
          59233 => x"00", -- $0e761
          59234 => x"00", -- $0e762
          59235 => x"00", -- $0e763
          59236 => x"00", -- $0e764
          59237 => x"00", -- $0e765
          59238 => x"00", -- $0e766
          59239 => x"00", -- $0e767
          59240 => x"00", -- $0e768
          59241 => x"00", -- $0e769
          59242 => x"00", -- $0e76a
          59243 => x"00", -- $0e76b
          59244 => x"00", -- $0e76c
          59245 => x"00", -- $0e76d
          59246 => x"00", -- $0e76e
          59247 => x"00", -- $0e76f
          59248 => x"00", -- $0e770
          59249 => x"00", -- $0e771
          59250 => x"00", -- $0e772
          59251 => x"00", -- $0e773
          59252 => x"00", -- $0e774
          59253 => x"00", -- $0e775
          59254 => x"00", -- $0e776
          59255 => x"00", -- $0e777
          59256 => x"00", -- $0e778
          59257 => x"00", -- $0e779
          59258 => x"00", -- $0e77a
          59259 => x"00", -- $0e77b
          59260 => x"00", -- $0e77c
          59261 => x"00", -- $0e77d
          59262 => x"00", -- $0e77e
          59263 => x"00", -- $0e77f
          59264 => x"00", -- $0e780
          59265 => x"00", -- $0e781
          59266 => x"00", -- $0e782
          59267 => x"00", -- $0e783
          59268 => x"00", -- $0e784
          59269 => x"00", -- $0e785
          59270 => x"00", -- $0e786
          59271 => x"00", -- $0e787
          59272 => x"00", -- $0e788
          59273 => x"00", -- $0e789
          59274 => x"00", -- $0e78a
          59275 => x"00", -- $0e78b
          59276 => x"00", -- $0e78c
          59277 => x"00", -- $0e78d
          59278 => x"00", -- $0e78e
          59279 => x"00", -- $0e78f
          59280 => x"00", -- $0e790
          59281 => x"00", -- $0e791
          59282 => x"00", -- $0e792
          59283 => x"00", -- $0e793
          59284 => x"00", -- $0e794
          59285 => x"00", -- $0e795
          59286 => x"00", -- $0e796
          59287 => x"00", -- $0e797
          59288 => x"00", -- $0e798
          59289 => x"00", -- $0e799
          59290 => x"00", -- $0e79a
          59291 => x"00", -- $0e79b
          59292 => x"00", -- $0e79c
          59293 => x"00", -- $0e79d
          59294 => x"00", -- $0e79e
          59295 => x"00", -- $0e79f
          59296 => x"00", -- $0e7a0
          59297 => x"00", -- $0e7a1
          59298 => x"00", -- $0e7a2
          59299 => x"00", -- $0e7a3
          59300 => x"00", -- $0e7a4
          59301 => x"00", -- $0e7a5
          59302 => x"00", -- $0e7a6
          59303 => x"00", -- $0e7a7
          59304 => x"00", -- $0e7a8
          59305 => x"00", -- $0e7a9
          59306 => x"00", -- $0e7aa
          59307 => x"00", -- $0e7ab
          59308 => x"00", -- $0e7ac
          59309 => x"00", -- $0e7ad
          59310 => x"00", -- $0e7ae
          59311 => x"00", -- $0e7af
          59312 => x"00", -- $0e7b0
          59313 => x"00", -- $0e7b1
          59314 => x"00", -- $0e7b2
          59315 => x"00", -- $0e7b3
          59316 => x"00", -- $0e7b4
          59317 => x"00", -- $0e7b5
          59318 => x"00", -- $0e7b6
          59319 => x"00", -- $0e7b7
          59320 => x"00", -- $0e7b8
          59321 => x"00", -- $0e7b9
          59322 => x"00", -- $0e7ba
          59323 => x"00", -- $0e7bb
          59324 => x"00", -- $0e7bc
          59325 => x"00", -- $0e7bd
          59326 => x"00", -- $0e7be
          59327 => x"00", -- $0e7bf
          59328 => x"00", -- $0e7c0
          59329 => x"00", -- $0e7c1
          59330 => x"00", -- $0e7c2
          59331 => x"00", -- $0e7c3
          59332 => x"00", -- $0e7c4
          59333 => x"00", -- $0e7c5
          59334 => x"00", -- $0e7c6
          59335 => x"00", -- $0e7c7
          59336 => x"00", -- $0e7c8
          59337 => x"00", -- $0e7c9
          59338 => x"00", -- $0e7ca
          59339 => x"00", -- $0e7cb
          59340 => x"00", -- $0e7cc
          59341 => x"00", -- $0e7cd
          59342 => x"00", -- $0e7ce
          59343 => x"00", -- $0e7cf
          59344 => x"00", -- $0e7d0
          59345 => x"00", -- $0e7d1
          59346 => x"00", -- $0e7d2
          59347 => x"00", -- $0e7d3
          59348 => x"00", -- $0e7d4
          59349 => x"00", -- $0e7d5
          59350 => x"00", -- $0e7d6
          59351 => x"00", -- $0e7d7
          59352 => x"00", -- $0e7d8
          59353 => x"00", -- $0e7d9
          59354 => x"00", -- $0e7da
          59355 => x"00", -- $0e7db
          59356 => x"00", -- $0e7dc
          59357 => x"00", -- $0e7dd
          59358 => x"00", -- $0e7de
          59359 => x"00", -- $0e7df
          59360 => x"00", -- $0e7e0
          59361 => x"00", -- $0e7e1
          59362 => x"00", -- $0e7e2
          59363 => x"00", -- $0e7e3
          59364 => x"00", -- $0e7e4
          59365 => x"00", -- $0e7e5
          59366 => x"00", -- $0e7e6
          59367 => x"00", -- $0e7e7
          59368 => x"00", -- $0e7e8
          59369 => x"00", -- $0e7e9
          59370 => x"00", -- $0e7ea
          59371 => x"00", -- $0e7eb
          59372 => x"00", -- $0e7ec
          59373 => x"00", -- $0e7ed
          59374 => x"00", -- $0e7ee
          59375 => x"00", -- $0e7ef
          59376 => x"00", -- $0e7f0
          59377 => x"00", -- $0e7f1
          59378 => x"00", -- $0e7f2
          59379 => x"00", -- $0e7f3
          59380 => x"00", -- $0e7f4
          59381 => x"00", -- $0e7f5
          59382 => x"00", -- $0e7f6
          59383 => x"00", -- $0e7f7
          59384 => x"00", -- $0e7f8
          59385 => x"00", -- $0e7f9
          59386 => x"00", -- $0e7fa
          59387 => x"00", -- $0e7fb
          59388 => x"00", -- $0e7fc
          59389 => x"00", -- $0e7fd
          59390 => x"00", -- $0e7fe
          59391 => x"00", -- $0e7ff
          59392 => x"00", -- $0e800
          59393 => x"00", -- $0e801
          59394 => x"00", -- $0e802
          59395 => x"00", -- $0e803
          59396 => x"00", -- $0e804
          59397 => x"00", -- $0e805
          59398 => x"00", -- $0e806
          59399 => x"00", -- $0e807
          59400 => x"00", -- $0e808
          59401 => x"00", -- $0e809
          59402 => x"00", -- $0e80a
          59403 => x"00", -- $0e80b
          59404 => x"00", -- $0e80c
          59405 => x"00", -- $0e80d
          59406 => x"00", -- $0e80e
          59407 => x"00", -- $0e80f
          59408 => x"00", -- $0e810
          59409 => x"00", -- $0e811
          59410 => x"00", -- $0e812
          59411 => x"00", -- $0e813
          59412 => x"00", -- $0e814
          59413 => x"00", -- $0e815
          59414 => x"00", -- $0e816
          59415 => x"00", -- $0e817
          59416 => x"00", -- $0e818
          59417 => x"00", -- $0e819
          59418 => x"00", -- $0e81a
          59419 => x"00", -- $0e81b
          59420 => x"00", -- $0e81c
          59421 => x"00", -- $0e81d
          59422 => x"00", -- $0e81e
          59423 => x"00", -- $0e81f
          59424 => x"00", -- $0e820
          59425 => x"00", -- $0e821
          59426 => x"00", -- $0e822
          59427 => x"00", -- $0e823
          59428 => x"00", -- $0e824
          59429 => x"00", -- $0e825
          59430 => x"00", -- $0e826
          59431 => x"00", -- $0e827
          59432 => x"00", -- $0e828
          59433 => x"00", -- $0e829
          59434 => x"00", -- $0e82a
          59435 => x"00", -- $0e82b
          59436 => x"00", -- $0e82c
          59437 => x"00", -- $0e82d
          59438 => x"00", -- $0e82e
          59439 => x"00", -- $0e82f
          59440 => x"00", -- $0e830
          59441 => x"00", -- $0e831
          59442 => x"00", -- $0e832
          59443 => x"00", -- $0e833
          59444 => x"00", -- $0e834
          59445 => x"00", -- $0e835
          59446 => x"00", -- $0e836
          59447 => x"00", -- $0e837
          59448 => x"00", -- $0e838
          59449 => x"00", -- $0e839
          59450 => x"00", -- $0e83a
          59451 => x"00", -- $0e83b
          59452 => x"00", -- $0e83c
          59453 => x"00", -- $0e83d
          59454 => x"00", -- $0e83e
          59455 => x"00", -- $0e83f
          59456 => x"00", -- $0e840
          59457 => x"00", -- $0e841
          59458 => x"00", -- $0e842
          59459 => x"00", -- $0e843
          59460 => x"00", -- $0e844
          59461 => x"00", -- $0e845
          59462 => x"00", -- $0e846
          59463 => x"00", -- $0e847
          59464 => x"00", -- $0e848
          59465 => x"00", -- $0e849
          59466 => x"00", -- $0e84a
          59467 => x"00", -- $0e84b
          59468 => x"00", -- $0e84c
          59469 => x"00", -- $0e84d
          59470 => x"00", -- $0e84e
          59471 => x"00", -- $0e84f
          59472 => x"00", -- $0e850
          59473 => x"00", -- $0e851
          59474 => x"00", -- $0e852
          59475 => x"00", -- $0e853
          59476 => x"00", -- $0e854
          59477 => x"00", -- $0e855
          59478 => x"00", -- $0e856
          59479 => x"00", -- $0e857
          59480 => x"00", -- $0e858
          59481 => x"00", -- $0e859
          59482 => x"00", -- $0e85a
          59483 => x"00", -- $0e85b
          59484 => x"00", -- $0e85c
          59485 => x"00", -- $0e85d
          59486 => x"00", -- $0e85e
          59487 => x"00", -- $0e85f
          59488 => x"00", -- $0e860
          59489 => x"00", -- $0e861
          59490 => x"00", -- $0e862
          59491 => x"00", -- $0e863
          59492 => x"00", -- $0e864
          59493 => x"00", -- $0e865
          59494 => x"00", -- $0e866
          59495 => x"00", -- $0e867
          59496 => x"00", -- $0e868
          59497 => x"00", -- $0e869
          59498 => x"00", -- $0e86a
          59499 => x"00", -- $0e86b
          59500 => x"00", -- $0e86c
          59501 => x"00", -- $0e86d
          59502 => x"00", -- $0e86e
          59503 => x"00", -- $0e86f
          59504 => x"00", -- $0e870
          59505 => x"00", -- $0e871
          59506 => x"00", -- $0e872
          59507 => x"00", -- $0e873
          59508 => x"00", -- $0e874
          59509 => x"00", -- $0e875
          59510 => x"00", -- $0e876
          59511 => x"00", -- $0e877
          59512 => x"00", -- $0e878
          59513 => x"00", -- $0e879
          59514 => x"00", -- $0e87a
          59515 => x"00", -- $0e87b
          59516 => x"00", -- $0e87c
          59517 => x"00", -- $0e87d
          59518 => x"00", -- $0e87e
          59519 => x"00", -- $0e87f
          59520 => x"00", -- $0e880
          59521 => x"00", -- $0e881
          59522 => x"00", -- $0e882
          59523 => x"00", -- $0e883
          59524 => x"00", -- $0e884
          59525 => x"00", -- $0e885
          59526 => x"00", -- $0e886
          59527 => x"00", -- $0e887
          59528 => x"00", -- $0e888
          59529 => x"00", -- $0e889
          59530 => x"00", -- $0e88a
          59531 => x"00", -- $0e88b
          59532 => x"00", -- $0e88c
          59533 => x"00", -- $0e88d
          59534 => x"00", -- $0e88e
          59535 => x"00", -- $0e88f
          59536 => x"00", -- $0e890
          59537 => x"00", -- $0e891
          59538 => x"00", -- $0e892
          59539 => x"00", -- $0e893
          59540 => x"00", -- $0e894
          59541 => x"00", -- $0e895
          59542 => x"00", -- $0e896
          59543 => x"00", -- $0e897
          59544 => x"00", -- $0e898
          59545 => x"00", -- $0e899
          59546 => x"00", -- $0e89a
          59547 => x"00", -- $0e89b
          59548 => x"00", -- $0e89c
          59549 => x"00", -- $0e89d
          59550 => x"00", -- $0e89e
          59551 => x"00", -- $0e89f
          59552 => x"00", -- $0e8a0
          59553 => x"00", -- $0e8a1
          59554 => x"00", -- $0e8a2
          59555 => x"00", -- $0e8a3
          59556 => x"00", -- $0e8a4
          59557 => x"00", -- $0e8a5
          59558 => x"00", -- $0e8a6
          59559 => x"00", -- $0e8a7
          59560 => x"00", -- $0e8a8
          59561 => x"00", -- $0e8a9
          59562 => x"00", -- $0e8aa
          59563 => x"00", -- $0e8ab
          59564 => x"00", -- $0e8ac
          59565 => x"00", -- $0e8ad
          59566 => x"00", -- $0e8ae
          59567 => x"00", -- $0e8af
          59568 => x"00", -- $0e8b0
          59569 => x"00", -- $0e8b1
          59570 => x"00", -- $0e8b2
          59571 => x"00", -- $0e8b3
          59572 => x"00", -- $0e8b4
          59573 => x"00", -- $0e8b5
          59574 => x"00", -- $0e8b6
          59575 => x"00", -- $0e8b7
          59576 => x"00", -- $0e8b8
          59577 => x"00", -- $0e8b9
          59578 => x"00", -- $0e8ba
          59579 => x"00", -- $0e8bb
          59580 => x"00", -- $0e8bc
          59581 => x"00", -- $0e8bd
          59582 => x"00", -- $0e8be
          59583 => x"00", -- $0e8bf
          59584 => x"00", -- $0e8c0
          59585 => x"00", -- $0e8c1
          59586 => x"00", -- $0e8c2
          59587 => x"00", -- $0e8c3
          59588 => x"00", -- $0e8c4
          59589 => x"00", -- $0e8c5
          59590 => x"00", -- $0e8c6
          59591 => x"00", -- $0e8c7
          59592 => x"00", -- $0e8c8
          59593 => x"00", -- $0e8c9
          59594 => x"00", -- $0e8ca
          59595 => x"00", -- $0e8cb
          59596 => x"00", -- $0e8cc
          59597 => x"00", -- $0e8cd
          59598 => x"00", -- $0e8ce
          59599 => x"00", -- $0e8cf
          59600 => x"00", -- $0e8d0
          59601 => x"00", -- $0e8d1
          59602 => x"00", -- $0e8d2
          59603 => x"00", -- $0e8d3
          59604 => x"00", -- $0e8d4
          59605 => x"00", -- $0e8d5
          59606 => x"00", -- $0e8d6
          59607 => x"00", -- $0e8d7
          59608 => x"00", -- $0e8d8
          59609 => x"00", -- $0e8d9
          59610 => x"00", -- $0e8da
          59611 => x"00", -- $0e8db
          59612 => x"00", -- $0e8dc
          59613 => x"00", -- $0e8dd
          59614 => x"00", -- $0e8de
          59615 => x"00", -- $0e8df
          59616 => x"00", -- $0e8e0
          59617 => x"00", -- $0e8e1
          59618 => x"00", -- $0e8e2
          59619 => x"00", -- $0e8e3
          59620 => x"00", -- $0e8e4
          59621 => x"00", -- $0e8e5
          59622 => x"00", -- $0e8e6
          59623 => x"00", -- $0e8e7
          59624 => x"00", -- $0e8e8
          59625 => x"00", -- $0e8e9
          59626 => x"00", -- $0e8ea
          59627 => x"00", -- $0e8eb
          59628 => x"00", -- $0e8ec
          59629 => x"00", -- $0e8ed
          59630 => x"00", -- $0e8ee
          59631 => x"00", -- $0e8ef
          59632 => x"00", -- $0e8f0
          59633 => x"00", -- $0e8f1
          59634 => x"00", -- $0e8f2
          59635 => x"00", -- $0e8f3
          59636 => x"00", -- $0e8f4
          59637 => x"00", -- $0e8f5
          59638 => x"00", -- $0e8f6
          59639 => x"00", -- $0e8f7
          59640 => x"00", -- $0e8f8
          59641 => x"00", -- $0e8f9
          59642 => x"00", -- $0e8fa
          59643 => x"00", -- $0e8fb
          59644 => x"00", -- $0e8fc
          59645 => x"00", -- $0e8fd
          59646 => x"00", -- $0e8fe
          59647 => x"00", -- $0e8ff
          59648 => x"00", -- $0e900
          59649 => x"00", -- $0e901
          59650 => x"00", -- $0e902
          59651 => x"00", -- $0e903
          59652 => x"00", -- $0e904
          59653 => x"00", -- $0e905
          59654 => x"00", -- $0e906
          59655 => x"00", -- $0e907
          59656 => x"00", -- $0e908
          59657 => x"00", -- $0e909
          59658 => x"00", -- $0e90a
          59659 => x"00", -- $0e90b
          59660 => x"00", -- $0e90c
          59661 => x"00", -- $0e90d
          59662 => x"00", -- $0e90e
          59663 => x"00", -- $0e90f
          59664 => x"00", -- $0e910
          59665 => x"00", -- $0e911
          59666 => x"00", -- $0e912
          59667 => x"00", -- $0e913
          59668 => x"00", -- $0e914
          59669 => x"00", -- $0e915
          59670 => x"00", -- $0e916
          59671 => x"00", -- $0e917
          59672 => x"00", -- $0e918
          59673 => x"00", -- $0e919
          59674 => x"00", -- $0e91a
          59675 => x"00", -- $0e91b
          59676 => x"00", -- $0e91c
          59677 => x"00", -- $0e91d
          59678 => x"00", -- $0e91e
          59679 => x"00", -- $0e91f
          59680 => x"00", -- $0e920
          59681 => x"00", -- $0e921
          59682 => x"00", -- $0e922
          59683 => x"00", -- $0e923
          59684 => x"00", -- $0e924
          59685 => x"00", -- $0e925
          59686 => x"00", -- $0e926
          59687 => x"00", -- $0e927
          59688 => x"00", -- $0e928
          59689 => x"00", -- $0e929
          59690 => x"00", -- $0e92a
          59691 => x"00", -- $0e92b
          59692 => x"00", -- $0e92c
          59693 => x"00", -- $0e92d
          59694 => x"00", -- $0e92e
          59695 => x"00", -- $0e92f
          59696 => x"00", -- $0e930
          59697 => x"00", -- $0e931
          59698 => x"00", -- $0e932
          59699 => x"00", -- $0e933
          59700 => x"00", -- $0e934
          59701 => x"00", -- $0e935
          59702 => x"00", -- $0e936
          59703 => x"00", -- $0e937
          59704 => x"00", -- $0e938
          59705 => x"00", -- $0e939
          59706 => x"00", -- $0e93a
          59707 => x"00", -- $0e93b
          59708 => x"00", -- $0e93c
          59709 => x"00", -- $0e93d
          59710 => x"00", -- $0e93e
          59711 => x"00", -- $0e93f
          59712 => x"00", -- $0e940
          59713 => x"00", -- $0e941
          59714 => x"00", -- $0e942
          59715 => x"00", -- $0e943
          59716 => x"00", -- $0e944
          59717 => x"00", -- $0e945
          59718 => x"00", -- $0e946
          59719 => x"00", -- $0e947
          59720 => x"00", -- $0e948
          59721 => x"00", -- $0e949
          59722 => x"00", -- $0e94a
          59723 => x"00", -- $0e94b
          59724 => x"00", -- $0e94c
          59725 => x"00", -- $0e94d
          59726 => x"00", -- $0e94e
          59727 => x"00", -- $0e94f
          59728 => x"00", -- $0e950
          59729 => x"00", -- $0e951
          59730 => x"00", -- $0e952
          59731 => x"00", -- $0e953
          59732 => x"00", -- $0e954
          59733 => x"00", -- $0e955
          59734 => x"00", -- $0e956
          59735 => x"00", -- $0e957
          59736 => x"00", -- $0e958
          59737 => x"00", -- $0e959
          59738 => x"00", -- $0e95a
          59739 => x"00", -- $0e95b
          59740 => x"00", -- $0e95c
          59741 => x"00", -- $0e95d
          59742 => x"00", -- $0e95e
          59743 => x"00", -- $0e95f
          59744 => x"00", -- $0e960
          59745 => x"00", -- $0e961
          59746 => x"00", -- $0e962
          59747 => x"00", -- $0e963
          59748 => x"00", -- $0e964
          59749 => x"00", -- $0e965
          59750 => x"00", -- $0e966
          59751 => x"00", -- $0e967
          59752 => x"00", -- $0e968
          59753 => x"00", -- $0e969
          59754 => x"00", -- $0e96a
          59755 => x"00", -- $0e96b
          59756 => x"00", -- $0e96c
          59757 => x"00", -- $0e96d
          59758 => x"00", -- $0e96e
          59759 => x"00", -- $0e96f
          59760 => x"00", -- $0e970
          59761 => x"00", -- $0e971
          59762 => x"00", -- $0e972
          59763 => x"00", -- $0e973
          59764 => x"00", -- $0e974
          59765 => x"00", -- $0e975
          59766 => x"00", -- $0e976
          59767 => x"00", -- $0e977
          59768 => x"00", -- $0e978
          59769 => x"00", -- $0e979
          59770 => x"00", -- $0e97a
          59771 => x"00", -- $0e97b
          59772 => x"00", -- $0e97c
          59773 => x"00", -- $0e97d
          59774 => x"00", -- $0e97e
          59775 => x"00", -- $0e97f
          59776 => x"00", -- $0e980
          59777 => x"00", -- $0e981
          59778 => x"00", -- $0e982
          59779 => x"00", -- $0e983
          59780 => x"00", -- $0e984
          59781 => x"00", -- $0e985
          59782 => x"00", -- $0e986
          59783 => x"00", -- $0e987
          59784 => x"00", -- $0e988
          59785 => x"00", -- $0e989
          59786 => x"00", -- $0e98a
          59787 => x"00", -- $0e98b
          59788 => x"00", -- $0e98c
          59789 => x"00", -- $0e98d
          59790 => x"00", -- $0e98e
          59791 => x"00", -- $0e98f
          59792 => x"00", -- $0e990
          59793 => x"00", -- $0e991
          59794 => x"00", -- $0e992
          59795 => x"00", -- $0e993
          59796 => x"00", -- $0e994
          59797 => x"00", -- $0e995
          59798 => x"00", -- $0e996
          59799 => x"00", -- $0e997
          59800 => x"00", -- $0e998
          59801 => x"00", -- $0e999
          59802 => x"00", -- $0e99a
          59803 => x"00", -- $0e99b
          59804 => x"00", -- $0e99c
          59805 => x"00", -- $0e99d
          59806 => x"00", -- $0e99e
          59807 => x"00", -- $0e99f
          59808 => x"00", -- $0e9a0
          59809 => x"00", -- $0e9a1
          59810 => x"00", -- $0e9a2
          59811 => x"00", -- $0e9a3
          59812 => x"00", -- $0e9a4
          59813 => x"00", -- $0e9a5
          59814 => x"00", -- $0e9a6
          59815 => x"00", -- $0e9a7
          59816 => x"00", -- $0e9a8
          59817 => x"00", -- $0e9a9
          59818 => x"00", -- $0e9aa
          59819 => x"00", -- $0e9ab
          59820 => x"00", -- $0e9ac
          59821 => x"00", -- $0e9ad
          59822 => x"00", -- $0e9ae
          59823 => x"00", -- $0e9af
          59824 => x"00", -- $0e9b0
          59825 => x"00", -- $0e9b1
          59826 => x"00", -- $0e9b2
          59827 => x"00", -- $0e9b3
          59828 => x"00", -- $0e9b4
          59829 => x"00", -- $0e9b5
          59830 => x"00", -- $0e9b6
          59831 => x"00", -- $0e9b7
          59832 => x"00", -- $0e9b8
          59833 => x"00", -- $0e9b9
          59834 => x"00", -- $0e9ba
          59835 => x"00", -- $0e9bb
          59836 => x"00", -- $0e9bc
          59837 => x"00", -- $0e9bd
          59838 => x"00", -- $0e9be
          59839 => x"00", -- $0e9bf
          59840 => x"00", -- $0e9c0
          59841 => x"00", -- $0e9c1
          59842 => x"00", -- $0e9c2
          59843 => x"00", -- $0e9c3
          59844 => x"00", -- $0e9c4
          59845 => x"00", -- $0e9c5
          59846 => x"00", -- $0e9c6
          59847 => x"00", -- $0e9c7
          59848 => x"00", -- $0e9c8
          59849 => x"00", -- $0e9c9
          59850 => x"00", -- $0e9ca
          59851 => x"00", -- $0e9cb
          59852 => x"00", -- $0e9cc
          59853 => x"00", -- $0e9cd
          59854 => x"00", -- $0e9ce
          59855 => x"00", -- $0e9cf
          59856 => x"00", -- $0e9d0
          59857 => x"00", -- $0e9d1
          59858 => x"00", -- $0e9d2
          59859 => x"00", -- $0e9d3
          59860 => x"00", -- $0e9d4
          59861 => x"00", -- $0e9d5
          59862 => x"00", -- $0e9d6
          59863 => x"00", -- $0e9d7
          59864 => x"00", -- $0e9d8
          59865 => x"00", -- $0e9d9
          59866 => x"00", -- $0e9da
          59867 => x"00", -- $0e9db
          59868 => x"00", -- $0e9dc
          59869 => x"00", -- $0e9dd
          59870 => x"00", -- $0e9de
          59871 => x"00", -- $0e9df
          59872 => x"00", -- $0e9e0
          59873 => x"00", -- $0e9e1
          59874 => x"00", -- $0e9e2
          59875 => x"00", -- $0e9e3
          59876 => x"00", -- $0e9e4
          59877 => x"00", -- $0e9e5
          59878 => x"00", -- $0e9e6
          59879 => x"00", -- $0e9e7
          59880 => x"00", -- $0e9e8
          59881 => x"00", -- $0e9e9
          59882 => x"00", -- $0e9ea
          59883 => x"00", -- $0e9eb
          59884 => x"00", -- $0e9ec
          59885 => x"00", -- $0e9ed
          59886 => x"00", -- $0e9ee
          59887 => x"00", -- $0e9ef
          59888 => x"00", -- $0e9f0
          59889 => x"00", -- $0e9f1
          59890 => x"00", -- $0e9f2
          59891 => x"00", -- $0e9f3
          59892 => x"00", -- $0e9f4
          59893 => x"00", -- $0e9f5
          59894 => x"00", -- $0e9f6
          59895 => x"00", -- $0e9f7
          59896 => x"00", -- $0e9f8
          59897 => x"00", -- $0e9f9
          59898 => x"00", -- $0e9fa
          59899 => x"00", -- $0e9fb
          59900 => x"00", -- $0e9fc
          59901 => x"00", -- $0e9fd
          59902 => x"00", -- $0e9fe
          59903 => x"00", -- $0e9ff
          59904 => x"00", -- $0ea00
          59905 => x"00", -- $0ea01
          59906 => x"00", -- $0ea02
          59907 => x"00", -- $0ea03
          59908 => x"00", -- $0ea04
          59909 => x"00", -- $0ea05
          59910 => x"00", -- $0ea06
          59911 => x"00", -- $0ea07
          59912 => x"00", -- $0ea08
          59913 => x"00", -- $0ea09
          59914 => x"00", -- $0ea0a
          59915 => x"00", -- $0ea0b
          59916 => x"00", -- $0ea0c
          59917 => x"00", -- $0ea0d
          59918 => x"00", -- $0ea0e
          59919 => x"00", -- $0ea0f
          59920 => x"00", -- $0ea10
          59921 => x"00", -- $0ea11
          59922 => x"00", -- $0ea12
          59923 => x"00", -- $0ea13
          59924 => x"00", -- $0ea14
          59925 => x"00", -- $0ea15
          59926 => x"00", -- $0ea16
          59927 => x"00", -- $0ea17
          59928 => x"00", -- $0ea18
          59929 => x"00", -- $0ea19
          59930 => x"00", -- $0ea1a
          59931 => x"00", -- $0ea1b
          59932 => x"00", -- $0ea1c
          59933 => x"00", -- $0ea1d
          59934 => x"00", -- $0ea1e
          59935 => x"00", -- $0ea1f
          59936 => x"00", -- $0ea20
          59937 => x"00", -- $0ea21
          59938 => x"00", -- $0ea22
          59939 => x"00", -- $0ea23
          59940 => x"00", -- $0ea24
          59941 => x"00", -- $0ea25
          59942 => x"00", -- $0ea26
          59943 => x"00", -- $0ea27
          59944 => x"00", -- $0ea28
          59945 => x"00", -- $0ea29
          59946 => x"00", -- $0ea2a
          59947 => x"00", -- $0ea2b
          59948 => x"00", -- $0ea2c
          59949 => x"00", -- $0ea2d
          59950 => x"00", -- $0ea2e
          59951 => x"00", -- $0ea2f
          59952 => x"00", -- $0ea30
          59953 => x"00", -- $0ea31
          59954 => x"00", -- $0ea32
          59955 => x"00", -- $0ea33
          59956 => x"00", -- $0ea34
          59957 => x"00", -- $0ea35
          59958 => x"00", -- $0ea36
          59959 => x"00", -- $0ea37
          59960 => x"00", -- $0ea38
          59961 => x"00", -- $0ea39
          59962 => x"00", -- $0ea3a
          59963 => x"00", -- $0ea3b
          59964 => x"00", -- $0ea3c
          59965 => x"00", -- $0ea3d
          59966 => x"00", -- $0ea3e
          59967 => x"00", -- $0ea3f
          59968 => x"00", -- $0ea40
          59969 => x"00", -- $0ea41
          59970 => x"00", -- $0ea42
          59971 => x"00", -- $0ea43
          59972 => x"00", -- $0ea44
          59973 => x"00", -- $0ea45
          59974 => x"00", -- $0ea46
          59975 => x"00", -- $0ea47
          59976 => x"00", -- $0ea48
          59977 => x"00", -- $0ea49
          59978 => x"00", -- $0ea4a
          59979 => x"00", -- $0ea4b
          59980 => x"00", -- $0ea4c
          59981 => x"00", -- $0ea4d
          59982 => x"00", -- $0ea4e
          59983 => x"00", -- $0ea4f
          59984 => x"00", -- $0ea50
          59985 => x"00", -- $0ea51
          59986 => x"00", -- $0ea52
          59987 => x"00", -- $0ea53
          59988 => x"00", -- $0ea54
          59989 => x"00", -- $0ea55
          59990 => x"00", -- $0ea56
          59991 => x"00", -- $0ea57
          59992 => x"00", -- $0ea58
          59993 => x"00", -- $0ea59
          59994 => x"00", -- $0ea5a
          59995 => x"00", -- $0ea5b
          59996 => x"00", -- $0ea5c
          59997 => x"00", -- $0ea5d
          59998 => x"00", -- $0ea5e
          59999 => x"00", -- $0ea5f
          60000 => x"00", -- $0ea60
          60001 => x"00", -- $0ea61
          60002 => x"00", -- $0ea62
          60003 => x"00", -- $0ea63
          60004 => x"00", -- $0ea64
          60005 => x"00", -- $0ea65
          60006 => x"00", -- $0ea66
          60007 => x"00", -- $0ea67
          60008 => x"00", -- $0ea68
          60009 => x"00", -- $0ea69
          60010 => x"00", -- $0ea6a
          60011 => x"00", -- $0ea6b
          60012 => x"00", -- $0ea6c
          60013 => x"00", -- $0ea6d
          60014 => x"00", -- $0ea6e
          60015 => x"00", -- $0ea6f
          60016 => x"00", -- $0ea70
          60017 => x"00", -- $0ea71
          60018 => x"00", -- $0ea72
          60019 => x"00", -- $0ea73
          60020 => x"00", -- $0ea74
          60021 => x"00", -- $0ea75
          60022 => x"00", -- $0ea76
          60023 => x"00", -- $0ea77
          60024 => x"00", -- $0ea78
          60025 => x"00", -- $0ea79
          60026 => x"00", -- $0ea7a
          60027 => x"00", -- $0ea7b
          60028 => x"00", -- $0ea7c
          60029 => x"00", -- $0ea7d
          60030 => x"00", -- $0ea7e
          60031 => x"00", -- $0ea7f
          60032 => x"00", -- $0ea80
          60033 => x"00", -- $0ea81
          60034 => x"00", -- $0ea82
          60035 => x"00", -- $0ea83
          60036 => x"00", -- $0ea84
          60037 => x"00", -- $0ea85
          60038 => x"00", -- $0ea86
          60039 => x"00", -- $0ea87
          60040 => x"00", -- $0ea88
          60041 => x"00", -- $0ea89
          60042 => x"00", -- $0ea8a
          60043 => x"00", -- $0ea8b
          60044 => x"00", -- $0ea8c
          60045 => x"00", -- $0ea8d
          60046 => x"00", -- $0ea8e
          60047 => x"00", -- $0ea8f
          60048 => x"00", -- $0ea90
          60049 => x"00", -- $0ea91
          60050 => x"00", -- $0ea92
          60051 => x"00", -- $0ea93
          60052 => x"00", -- $0ea94
          60053 => x"00", -- $0ea95
          60054 => x"00", -- $0ea96
          60055 => x"00", -- $0ea97
          60056 => x"00", -- $0ea98
          60057 => x"00", -- $0ea99
          60058 => x"00", -- $0ea9a
          60059 => x"00", -- $0ea9b
          60060 => x"00", -- $0ea9c
          60061 => x"00", -- $0ea9d
          60062 => x"00", -- $0ea9e
          60063 => x"00", -- $0ea9f
          60064 => x"00", -- $0eaa0
          60065 => x"00", -- $0eaa1
          60066 => x"00", -- $0eaa2
          60067 => x"00", -- $0eaa3
          60068 => x"00", -- $0eaa4
          60069 => x"00", -- $0eaa5
          60070 => x"00", -- $0eaa6
          60071 => x"00", -- $0eaa7
          60072 => x"00", -- $0eaa8
          60073 => x"00", -- $0eaa9
          60074 => x"00", -- $0eaaa
          60075 => x"00", -- $0eaab
          60076 => x"00", -- $0eaac
          60077 => x"00", -- $0eaad
          60078 => x"00", -- $0eaae
          60079 => x"00", -- $0eaaf
          60080 => x"00", -- $0eab0
          60081 => x"00", -- $0eab1
          60082 => x"00", -- $0eab2
          60083 => x"00", -- $0eab3
          60084 => x"00", -- $0eab4
          60085 => x"00", -- $0eab5
          60086 => x"00", -- $0eab6
          60087 => x"00", -- $0eab7
          60088 => x"00", -- $0eab8
          60089 => x"00", -- $0eab9
          60090 => x"00", -- $0eaba
          60091 => x"00", -- $0eabb
          60092 => x"00", -- $0eabc
          60093 => x"00", -- $0eabd
          60094 => x"00", -- $0eabe
          60095 => x"00", -- $0eabf
          60096 => x"00", -- $0eac0
          60097 => x"00", -- $0eac1
          60098 => x"00", -- $0eac2
          60099 => x"00", -- $0eac3
          60100 => x"00", -- $0eac4
          60101 => x"00", -- $0eac5
          60102 => x"00", -- $0eac6
          60103 => x"00", -- $0eac7
          60104 => x"00", -- $0eac8
          60105 => x"00", -- $0eac9
          60106 => x"00", -- $0eaca
          60107 => x"00", -- $0eacb
          60108 => x"00", -- $0eacc
          60109 => x"00", -- $0eacd
          60110 => x"00", -- $0eace
          60111 => x"00", -- $0eacf
          60112 => x"00", -- $0ead0
          60113 => x"00", -- $0ead1
          60114 => x"00", -- $0ead2
          60115 => x"00", -- $0ead3
          60116 => x"00", -- $0ead4
          60117 => x"00", -- $0ead5
          60118 => x"00", -- $0ead6
          60119 => x"00", -- $0ead7
          60120 => x"00", -- $0ead8
          60121 => x"00", -- $0ead9
          60122 => x"00", -- $0eada
          60123 => x"00", -- $0eadb
          60124 => x"00", -- $0eadc
          60125 => x"00", -- $0eadd
          60126 => x"00", -- $0eade
          60127 => x"00", -- $0eadf
          60128 => x"00", -- $0eae0
          60129 => x"00", -- $0eae1
          60130 => x"00", -- $0eae2
          60131 => x"00", -- $0eae3
          60132 => x"00", -- $0eae4
          60133 => x"00", -- $0eae5
          60134 => x"00", -- $0eae6
          60135 => x"00", -- $0eae7
          60136 => x"00", -- $0eae8
          60137 => x"00", -- $0eae9
          60138 => x"00", -- $0eaea
          60139 => x"00", -- $0eaeb
          60140 => x"00", -- $0eaec
          60141 => x"00", -- $0eaed
          60142 => x"00", -- $0eaee
          60143 => x"00", -- $0eaef
          60144 => x"00", -- $0eaf0
          60145 => x"00", -- $0eaf1
          60146 => x"00", -- $0eaf2
          60147 => x"00", -- $0eaf3
          60148 => x"00", -- $0eaf4
          60149 => x"00", -- $0eaf5
          60150 => x"00", -- $0eaf6
          60151 => x"00", -- $0eaf7
          60152 => x"00", -- $0eaf8
          60153 => x"00", -- $0eaf9
          60154 => x"00", -- $0eafa
          60155 => x"00", -- $0eafb
          60156 => x"00", -- $0eafc
          60157 => x"00", -- $0eafd
          60158 => x"00", -- $0eafe
          60159 => x"00", -- $0eaff
          60160 => x"00", -- $0eb00
          60161 => x"00", -- $0eb01
          60162 => x"00", -- $0eb02
          60163 => x"00", -- $0eb03
          60164 => x"00", -- $0eb04
          60165 => x"00", -- $0eb05
          60166 => x"00", -- $0eb06
          60167 => x"00", -- $0eb07
          60168 => x"00", -- $0eb08
          60169 => x"00", -- $0eb09
          60170 => x"00", -- $0eb0a
          60171 => x"00", -- $0eb0b
          60172 => x"00", -- $0eb0c
          60173 => x"00", -- $0eb0d
          60174 => x"00", -- $0eb0e
          60175 => x"00", -- $0eb0f
          60176 => x"00", -- $0eb10
          60177 => x"00", -- $0eb11
          60178 => x"00", -- $0eb12
          60179 => x"00", -- $0eb13
          60180 => x"00", -- $0eb14
          60181 => x"00", -- $0eb15
          60182 => x"00", -- $0eb16
          60183 => x"00", -- $0eb17
          60184 => x"00", -- $0eb18
          60185 => x"00", -- $0eb19
          60186 => x"00", -- $0eb1a
          60187 => x"00", -- $0eb1b
          60188 => x"00", -- $0eb1c
          60189 => x"00", -- $0eb1d
          60190 => x"00", -- $0eb1e
          60191 => x"00", -- $0eb1f
          60192 => x"00", -- $0eb20
          60193 => x"00", -- $0eb21
          60194 => x"00", -- $0eb22
          60195 => x"00", -- $0eb23
          60196 => x"00", -- $0eb24
          60197 => x"00", -- $0eb25
          60198 => x"00", -- $0eb26
          60199 => x"00", -- $0eb27
          60200 => x"00", -- $0eb28
          60201 => x"00", -- $0eb29
          60202 => x"00", -- $0eb2a
          60203 => x"00", -- $0eb2b
          60204 => x"00", -- $0eb2c
          60205 => x"00", -- $0eb2d
          60206 => x"00", -- $0eb2e
          60207 => x"00", -- $0eb2f
          60208 => x"00", -- $0eb30
          60209 => x"00", -- $0eb31
          60210 => x"00", -- $0eb32
          60211 => x"00", -- $0eb33
          60212 => x"00", -- $0eb34
          60213 => x"00", -- $0eb35
          60214 => x"00", -- $0eb36
          60215 => x"00", -- $0eb37
          60216 => x"00", -- $0eb38
          60217 => x"00", -- $0eb39
          60218 => x"00", -- $0eb3a
          60219 => x"00", -- $0eb3b
          60220 => x"00", -- $0eb3c
          60221 => x"00", -- $0eb3d
          60222 => x"00", -- $0eb3e
          60223 => x"00", -- $0eb3f
          60224 => x"00", -- $0eb40
          60225 => x"00", -- $0eb41
          60226 => x"00", -- $0eb42
          60227 => x"00", -- $0eb43
          60228 => x"00", -- $0eb44
          60229 => x"00", -- $0eb45
          60230 => x"00", -- $0eb46
          60231 => x"00", -- $0eb47
          60232 => x"00", -- $0eb48
          60233 => x"00", -- $0eb49
          60234 => x"00", -- $0eb4a
          60235 => x"00", -- $0eb4b
          60236 => x"00", -- $0eb4c
          60237 => x"00", -- $0eb4d
          60238 => x"00", -- $0eb4e
          60239 => x"00", -- $0eb4f
          60240 => x"00", -- $0eb50
          60241 => x"00", -- $0eb51
          60242 => x"00", -- $0eb52
          60243 => x"00", -- $0eb53
          60244 => x"00", -- $0eb54
          60245 => x"00", -- $0eb55
          60246 => x"00", -- $0eb56
          60247 => x"00", -- $0eb57
          60248 => x"00", -- $0eb58
          60249 => x"00", -- $0eb59
          60250 => x"00", -- $0eb5a
          60251 => x"00", -- $0eb5b
          60252 => x"00", -- $0eb5c
          60253 => x"00", -- $0eb5d
          60254 => x"00", -- $0eb5e
          60255 => x"00", -- $0eb5f
          60256 => x"00", -- $0eb60
          60257 => x"00", -- $0eb61
          60258 => x"00", -- $0eb62
          60259 => x"00", -- $0eb63
          60260 => x"00", -- $0eb64
          60261 => x"00", -- $0eb65
          60262 => x"00", -- $0eb66
          60263 => x"00", -- $0eb67
          60264 => x"00", -- $0eb68
          60265 => x"00", -- $0eb69
          60266 => x"00", -- $0eb6a
          60267 => x"00", -- $0eb6b
          60268 => x"00", -- $0eb6c
          60269 => x"00", -- $0eb6d
          60270 => x"00", -- $0eb6e
          60271 => x"00", -- $0eb6f
          60272 => x"00", -- $0eb70
          60273 => x"00", -- $0eb71
          60274 => x"00", -- $0eb72
          60275 => x"00", -- $0eb73
          60276 => x"00", -- $0eb74
          60277 => x"00", -- $0eb75
          60278 => x"00", -- $0eb76
          60279 => x"00", -- $0eb77
          60280 => x"00", -- $0eb78
          60281 => x"00", -- $0eb79
          60282 => x"00", -- $0eb7a
          60283 => x"00", -- $0eb7b
          60284 => x"00", -- $0eb7c
          60285 => x"00", -- $0eb7d
          60286 => x"00", -- $0eb7e
          60287 => x"00", -- $0eb7f
          60288 => x"00", -- $0eb80
          60289 => x"00", -- $0eb81
          60290 => x"00", -- $0eb82
          60291 => x"00", -- $0eb83
          60292 => x"00", -- $0eb84
          60293 => x"00", -- $0eb85
          60294 => x"00", -- $0eb86
          60295 => x"00", -- $0eb87
          60296 => x"00", -- $0eb88
          60297 => x"00", -- $0eb89
          60298 => x"00", -- $0eb8a
          60299 => x"00", -- $0eb8b
          60300 => x"00", -- $0eb8c
          60301 => x"00", -- $0eb8d
          60302 => x"00", -- $0eb8e
          60303 => x"00", -- $0eb8f
          60304 => x"00", -- $0eb90
          60305 => x"00", -- $0eb91
          60306 => x"00", -- $0eb92
          60307 => x"00", -- $0eb93
          60308 => x"00", -- $0eb94
          60309 => x"00", -- $0eb95
          60310 => x"00", -- $0eb96
          60311 => x"00", -- $0eb97
          60312 => x"00", -- $0eb98
          60313 => x"00", -- $0eb99
          60314 => x"00", -- $0eb9a
          60315 => x"00", -- $0eb9b
          60316 => x"00", -- $0eb9c
          60317 => x"00", -- $0eb9d
          60318 => x"00", -- $0eb9e
          60319 => x"00", -- $0eb9f
          60320 => x"00", -- $0eba0
          60321 => x"00", -- $0eba1
          60322 => x"00", -- $0eba2
          60323 => x"00", -- $0eba3
          60324 => x"00", -- $0eba4
          60325 => x"00", -- $0eba5
          60326 => x"00", -- $0eba6
          60327 => x"00", -- $0eba7
          60328 => x"00", -- $0eba8
          60329 => x"00", -- $0eba9
          60330 => x"00", -- $0ebaa
          60331 => x"00", -- $0ebab
          60332 => x"00", -- $0ebac
          60333 => x"00", -- $0ebad
          60334 => x"00", -- $0ebae
          60335 => x"00", -- $0ebaf
          60336 => x"00", -- $0ebb0
          60337 => x"00", -- $0ebb1
          60338 => x"00", -- $0ebb2
          60339 => x"00", -- $0ebb3
          60340 => x"00", -- $0ebb4
          60341 => x"00", -- $0ebb5
          60342 => x"00", -- $0ebb6
          60343 => x"00", -- $0ebb7
          60344 => x"00", -- $0ebb8
          60345 => x"00", -- $0ebb9
          60346 => x"00", -- $0ebba
          60347 => x"00", -- $0ebbb
          60348 => x"00", -- $0ebbc
          60349 => x"00", -- $0ebbd
          60350 => x"00", -- $0ebbe
          60351 => x"00", -- $0ebbf
          60352 => x"00", -- $0ebc0
          60353 => x"00", -- $0ebc1
          60354 => x"00", -- $0ebc2
          60355 => x"00", -- $0ebc3
          60356 => x"00", -- $0ebc4
          60357 => x"00", -- $0ebc5
          60358 => x"00", -- $0ebc6
          60359 => x"00", -- $0ebc7
          60360 => x"00", -- $0ebc8
          60361 => x"00", -- $0ebc9
          60362 => x"00", -- $0ebca
          60363 => x"00", -- $0ebcb
          60364 => x"00", -- $0ebcc
          60365 => x"00", -- $0ebcd
          60366 => x"00", -- $0ebce
          60367 => x"00", -- $0ebcf
          60368 => x"00", -- $0ebd0
          60369 => x"00", -- $0ebd1
          60370 => x"00", -- $0ebd2
          60371 => x"00", -- $0ebd3
          60372 => x"00", -- $0ebd4
          60373 => x"00", -- $0ebd5
          60374 => x"00", -- $0ebd6
          60375 => x"00", -- $0ebd7
          60376 => x"00", -- $0ebd8
          60377 => x"00", -- $0ebd9
          60378 => x"00", -- $0ebda
          60379 => x"00", -- $0ebdb
          60380 => x"00", -- $0ebdc
          60381 => x"00", -- $0ebdd
          60382 => x"00", -- $0ebde
          60383 => x"00", -- $0ebdf
          60384 => x"00", -- $0ebe0
          60385 => x"00", -- $0ebe1
          60386 => x"00", -- $0ebe2
          60387 => x"00", -- $0ebe3
          60388 => x"00", -- $0ebe4
          60389 => x"00", -- $0ebe5
          60390 => x"00", -- $0ebe6
          60391 => x"00", -- $0ebe7
          60392 => x"00", -- $0ebe8
          60393 => x"00", -- $0ebe9
          60394 => x"00", -- $0ebea
          60395 => x"00", -- $0ebeb
          60396 => x"00", -- $0ebec
          60397 => x"00", -- $0ebed
          60398 => x"00", -- $0ebee
          60399 => x"00", -- $0ebef
          60400 => x"00", -- $0ebf0
          60401 => x"00", -- $0ebf1
          60402 => x"00", -- $0ebf2
          60403 => x"00", -- $0ebf3
          60404 => x"00", -- $0ebf4
          60405 => x"00", -- $0ebf5
          60406 => x"00", -- $0ebf6
          60407 => x"00", -- $0ebf7
          60408 => x"00", -- $0ebf8
          60409 => x"00", -- $0ebf9
          60410 => x"00", -- $0ebfa
          60411 => x"00", -- $0ebfb
          60412 => x"00", -- $0ebfc
          60413 => x"00", -- $0ebfd
          60414 => x"00", -- $0ebfe
          60415 => x"00", -- $0ebff
          60416 => x"00", -- $0ec00
          60417 => x"00", -- $0ec01
          60418 => x"00", -- $0ec02
          60419 => x"00", -- $0ec03
          60420 => x"00", -- $0ec04
          60421 => x"00", -- $0ec05
          60422 => x"00", -- $0ec06
          60423 => x"00", -- $0ec07
          60424 => x"00", -- $0ec08
          60425 => x"00", -- $0ec09
          60426 => x"00", -- $0ec0a
          60427 => x"00", -- $0ec0b
          60428 => x"00", -- $0ec0c
          60429 => x"00", -- $0ec0d
          60430 => x"00", -- $0ec0e
          60431 => x"00", -- $0ec0f
          60432 => x"00", -- $0ec10
          60433 => x"00", -- $0ec11
          60434 => x"00", -- $0ec12
          60435 => x"00", -- $0ec13
          60436 => x"00", -- $0ec14
          60437 => x"00", -- $0ec15
          60438 => x"00", -- $0ec16
          60439 => x"00", -- $0ec17
          60440 => x"00", -- $0ec18
          60441 => x"00", -- $0ec19
          60442 => x"00", -- $0ec1a
          60443 => x"00", -- $0ec1b
          60444 => x"00", -- $0ec1c
          60445 => x"00", -- $0ec1d
          60446 => x"00", -- $0ec1e
          60447 => x"00", -- $0ec1f
          60448 => x"00", -- $0ec20
          60449 => x"00", -- $0ec21
          60450 => x"00", -- $0ec22
          60451 => x"00", -- $0ec23
          60452 => x"00", -- $0ec24
          60453 => x"00", -- $0ec25
          60454 => x"00", -- $0ec26
          60455 => x"00", -- $0ec27
          60456 => x"00", -- $0ec28
          60457 => x"00", -- $0ec29
          60458 => x"00", -- $0ec2a
          60459 => x"00", -- $0ec2b
          60460 => x"00", -- $0ec2c
          60461 => x"00", -- $0ec2d
          60462 => x"00", -- $0ec2e
          60463 => x"00", -- $0ec2f
          60464 => x"00", -- $0ec30
          60465 => x"00", -- $0ec31
          60466 => x"00", -- $0ec32
          60467 => x"00", -- $0ec33
          60468 => x"00", -- $0ec34
          60469 => x"00", -- $0ec35
          60470 => x"00", -- $0ec36
          60471 => x"00", -- $0ec37
          60472 => x"00", -- $0ec38
          60473 => x"00", -- $0ec39
          60474 => x"00", -- $0ec3a
          60475 => x"00", -- $0ec3b
          60476 => x"00", -- $0ec3c
          60477 => x"00", -- $0ec3d
          60478 => x"00", -- $0ec3e
          60479 => x"00", -- $0ec3f
          60480 => x"00", -- $0ec40
          60481 => x"00", -- $0ec41
          60482 => x"00", -- $0ec42
          60483 => x"00", -- $0ec43
          60484 => x"00", -- $0ec44
          60485 => x"00", -- $0ec45
          60486 => x"00", -- $0ec46
          60487 => x"00", -- $0ec47
          60488 => x"00", -- $0ec48
          60489 => x"00", -- $0ec49
          60490 => x"00", -- $0ec4a
          60491 => x"00", -- $0ec4b
          60492 => x"00", -- $0ec4c
          60493 => x"00", -- $0ec4d
          60494 => x"00", -- $0ec4e
          60495 => x"00", -- $0ec4f
          60496 => x"00", -- $0ec50
          60497 => x"00", -- $0ec51
          60498 => x"00", -- $0ec52
          60499 => x"00", -- $0ec53
          60500 => x"00", -- $0ec54
          60501 => x"00", -- $0ec55
          60502 => x"00", -- $0ec56
          60503 => x"00", -- $0ec57
          60504 => x"00", -- $0ec58
          60505 => x"00", -- $0ec59
          60506 => x"00", -- $0ec5a
          60507 => x"00", -- $0ec5b
          60508 => x"00", -- $0ec5c
          60509 => x"00", -- $0ec5d
          60510 => x"00", -- $0ec5e
          60511 => x"00", -- $0ec5f
          60512 => x"00", -- $0ec60
          60513 => x"00", -- $0ec61
          60514 => x"00", -- $0ec62
          60515 => x"00", -- $0ec63
          60516 => x"00", -- $0ec64
          60517 => x"00", -- $0ec65
          60518 => x"00", -- $0ec66
          60519 => x"00", -- $0ec67
          60520 => x"00", -- $0ec68
          60521 => x"00", -- $0ec69
          60522 => x"00", -- $0ec6a
          60523 => x"00", -- $0ec6b
          60524 => x"00", -- $0ec6c
          60525 => x"00", -- $0ec6d
          60526 => x"00", -- $0ec6e
          60527 => x"00", -- $0ec6f
          60528 => x"00", -- $0ec70
          60529 => x"00", -- $0ec71
          60530 => x"00", -- $0ec72
          60531 => x"00", -- $0ec73
          60532 => x"00", -- $0ec74
          60533 => x"00", -- $0ec75
          60534 => x"00", -- $0ec76
          60535 => x"00", -- $0ec77
          60536 => x"00", -- $0ec78
          60537 => x"00", -- $0ec79
          60538 => x"00", -- $0ec7a
          60539 => x"00", -- $0ec7b
          60540 => x"00", -- $0ec7c
          60541 => x"00", -- $0ec7d
          60542 => x"00", -- $0ec7e
          60543 => x"00", -- $0ec7f
          60544 => x"00", -- $0ec80
          60545 => x"00", -- $0ec81
          60546 => x"00", -- $0ec82
          60547 => x"00", -- $0ec83
          60548 => x"00", -- $0ec84
          60549 => x"00", -- $0ec85
          60550 => x"00", -- $0ec86
          60551 => x"00", -- $0ec87
          60552 => x"00", -- $0ec88
          60553 => x"00", -- $0ec89
          60554 => x"00", -- $0ec8a
          60555 => x"00", -- $0ec8b
          60556 => x"00", -- $0ec8c
          60557 => x"00", -- $0ec8d
          60558 => x"00", -- $0ec8e
          60559 => x"00", -- $0ec8f
          60560 => x"00", -- $0ec90
          60561 => x"00", -- $0ec91
          60562 => x"00", -- $0ec92
          60563 => x"00", -- $0ec93
          60564 => x"00", -- $0ec94
          60565 => x"00", -- $0ec95
          60566 => x"00", -- $0ec96
          60567 => x"00", -- $0ec97
          60568 => x"00", -- $0ec98
          60569 => x"00", -- $0ec99
          60570 => x"00", -- $0ec9a
          60571 => x"00", -- $0ec9b
          60572 => x"00", -- $0ec9c
          60573 => x"00", -- $0ec9d
          60574 => x"00", -- $0ec9e
          60575 => x"00", -- $0ec9f
          60576 => x"00", -- $0eca0
          60577 => x"00", -- $0eca1
          60578 => x"00", -- $0eca2
          60579 => x"00", -- $0eca3
          60580 => x"00", -- $0eca4
          60581 => x"00", -- $0eca5
          60582 => x"00", -- $0eca6
          60583 => x"00", -- $0eca7
          60584 => x"00", -- $0eca8
          60585 => x"00", -- $0eca9
          60586 => x"00", -- $0ecaa
          60587 => x"00", -- $0ecab
          60588 => x"00", -- $0ecac
          60589 => x"00", -- $0ecad
          60590 => x"00", -- $0ecae
          60591 => x"00", -- $0ecaf
          60592 => x"00", -- $0ecb0
          60593 => x"00", -- $0ecb1
          60594 => x"00", -- $0ecb2
          60595 => x"00", -- $0ecb3
          60596 => x"00", -- $0ecb4
          60597 => x"00", -- $0ecb5
          60598 => x"00", -- $0ecb6
          60599 => x"00", -- $0ecb7
          60600 => x"00", -- $0ecb8
          60601 => x"00", -- $0ecb9
          60602 => x"00", -- $0ecba
          60603 => x"00", -- $0ecbb
          60604 => x"00", -- $0ecbc
          60605 => x"00", -- $0ecbd
          60606 => x"00", -- $0ecbe
          60607 => x"00", -- $0ecbf
          60608 => x"00", -- $0ecc0
          60609 => x"00", -- $0ecc1
          60610 => x"00", -- $0ecc2
          60611 => x"00", -- $0ecc3
          60612 => x"00", -- $0ecc4
          60613 => x"00", -- $0ecc5
          60614 => x"00", -- $0ecc6
          60615 => x"00", -- $0ecc7
          60616 => x"00", -- $0ecc8
          60617 => x"00", -- $0ecc9
          60618 => x"00", -- $0ecca
          60619 => x"00", -- $0eccb
          60620 => x"00", -- $0eccc
          60621 => x"00", -- $0eccd
          60622 => x"00", -- $0ecce
          60623 => x"00", -- $0eccf
          60624 => x"00", -- $0ecd0
          60625 => x"00", -- $0ecd1
          60626 => x"00", -- $0ecd2
          60627 => x"00", -- $0ecd3
          60628 => x"00", -- $0ecd4
          60629 => x"00", -- $0ecd5
          60630 => x"00", -- $0ecd6
          60631 => x"00", -- $0ecd7
          60632 => x"00", -- $0ecd8
          60633 => x"00", -- $0ecd9
          60634 => x"00", -- $0ecda
          60635 => x"00", -- $0ecdb
          60636 => x"00", -- $0ecdc
          60637 => x"00", -- $0ecdd
          60638 => x"00", -- $0ecde
          60639 => x"00", -- $0ecdf
          60640 => x"00", -- $0ece0
          60641 => x"00", -- $0ece1
          60642 => x"00", -- $0ece2
          60643 => x"00", -- $0ece3
          60644 => x"00", -- $0ece4
          60645 => x"00", -- $0ece5
          60646 => x"00", -- $0ece6
          60647 => x"00", -- $0ece7
          60648 => x"00", -- $0ece8
          60649 => x"00", -- $0ece9
          60650 => x"00", -- $0ecea
          60651 => x"00", -- $0eceb
          60652 => x"00", -- $0ecec
          60653 => x"00", -- $0eced
          60654 => x"00", -- $0ecee
          60655 => x"00", -- $0ecef
          60656 => x"00", -- $0ecf0
          60657 => x"00", -- $0ecf1
          60658 => x"00", -- $0ecf2
          60659 => x"00", -- $0ecf3
          60660 => x"00", -- $0ecf4
          60661 => x"00", -- $0ecf5
          60662 => x"00", -- $0ecf6
          60663 => x"00", -- $0ecf7
          60664 => x"00", -- $0ecf8
          60665 => x"00", -- $0ecf9
          60666 => x"00", -- $0ecfa
          60667 => x"00", -- $0ecfb
          60668 => x"00", -- $0ecfc
          60669 => x"00", -- $0ecfd
          60670 => x"00", -- $0ecfe
          60671 => x"00", -- $0ecff
          60672 => x"00", -- $0ed00
          60673 => x"00", -- $0ed01
          60674 => x"00", -- $0ed02
          60675 => x"00", -- $0ed03
          60676 => x"00", -- $0ed04
          60677 => x"00", -- $0ed05
          60678 => x"00", -- $0ed06
          60679 => x"00", -- $0ed07
          60680 => x"00", -- $0ed08
          60681 => x"00", -- $0ed09
          60682 => x"00", -- $0ed0a
          60683 => x"00", -- $0ed0b
          60684 => x"00", -- $0ed0c
          60685 => x"00", -- $0ed0d
          60686 => x"00", -- $0ed0e
          60687 => x"00", -- $0ed0f
          60688 => x"00", -- $0ed10
          60689 => x"00", -- $0ed11
          60690 => x"00", -- $0ed12
          60691 => x"00", -- $0ed13
          60692 => x"00", -- $0ed14
          60693 => x"00", -- $0ed15
          60694 => x"00", -- $0ed16
          60695 => x"00", -- $0ed17
          60696 => x"00", -- $0ed18
          60697 => x"00", -- $0ed19
          60698 => x"00", -- $0ed1a
          60699 => x"00", -- $0ed1b
          60700 => x"00", -- $0ed1c
          60701 => x"00", -- $0ed1d
          60702 => x"00", -- $0ed1e
          60703 => x"00", -- $0ed1f
          60704 => x"00", -- $0ed20
          60705 => x"00", -- $0ed21
          60706 => x"00", -- $0ed22
          60707 => x"00", -- $0ed23
          60708 => x"00", -- $0ed24
          60709 => x"00", -- $0ed25
          60710 => x"00", -- $0ed26
          60711 => x"00", -- $0ed27
          60712 => x"00", -- $0ed28
          60713 => x"00", -- $0ed29
          60714 => x"00", -- $0ed2a
          60715 => x"00", -- $0ed2b
          60716 => x"00", -- $0ed2c
          60717 => x"00", -- $0ed2d
          60718 => x"00", -- $0ed2e
          60719 => x"00", -- $0ed2f
          60720 => x"00", -- $0ed30
          60721 => x"00", -- $0ed31
          60722 => x"00", -- $0ed32
          60723 => x"00", -- $0ed33
          60724 => x"00", -- $0ed34
          60725 => x"00", -- $0ed35
          60726 => x"00", -- $0ed36
          60727 => x"00", -- $0ed37
          60728 => x"00", -- $0ed38
          60729 => x"00", -- $0ed39
          60730 => x"00", -- $0ed3a
          60731 => x"00", -- $0ed3b
          60732 => x"00", -- $0ed3c
          60733 => x"00", -- $0ed3d
          60734 => x"00", -- $0ed3e
          60735 => x"00", -- $0ed3f
          60736 => x"00", -- $0ed40
          60737 => x"00", -- $0ed41
          60738 => x"00", -- $0ed42
          60739 => x"00", -- $0ed43
          60740 => x"00", -- $0ed44
          60741 => x"00", -- $0ed45
          60742 => x"00", -- $0ed46
          60743 => x"00", -- $0ed47
          60744 => x"00", -- $0ed48
          60745 => x"00", -- $0ed49
          60746 => x"00", -- $0ed4a
          60747 => x"00", -- $0ed4b
          60748 => x"00", -- $0ed4c
          60749 => x"00", -- $0ed4d
          60750 => x"00", -- $0ed4e
          60751 => x"00", -- $0ed4f
          60752 => x"00", -- $0ed50
          60753 => x"00", -- $0ed51
          60754 => x"00", -- $0ed52
          60755 => x"00", -- $0ed53
          60756 => x"00", -- $0ed54
          60757 => x"00", -- $0ed55
          60758 => x"00", -- $0ed56
          60759 => x"00", -- $0ed57
          60760 => x"00", -- $0ed58
          60761 => x"00", -- $0ed59
          60762 => x"00", -- $0ed5a
          60763 => x"00", -- $0ed5b
          60764 => x"00", -- $0ed5c
          60765 => x"00", -- $0ed5d
          60766 => x"00", -- $0ed5e
          60767 => x"00", -- $0ed5f
          60768 => x"00", -- $0ed60
          60769 => x"00", -- $0ed61
          60770 => x"00", -- $0ed62
          60771 => x"00", -- $0ed63
          60772 => x"00", -- $0ed64
          60773 => x"00", -- $0ed65
          60774 => x"00", -- $0ed66
          60775 => x"00", -- $0ed67
          60776 => x"00", -- $0ed68
          60777 => x"00", -- $0ed69
          60778 => x"00", -- $0ed6a
          60779 => x"00", -- $0ed6b
          60780 => x"00", -- $0ed6c
          60781 => x"00", -- $0ed6d
          60782 => x"00", -- $0ed6e
          60783 => x"00", -- $0ed6f
          60784 => x"00", -- $0ed70
          60785 => x"00", -- $0ed71
          60786 => x"00", -- $0ed72
          60787 => x"00", -- $0ed73
          60788 => x"00", -- $0ed74
          60789 => x"00", -- $0ed75
          60790 => x"00", -- $0ed76
          60791 => x"00", -- $0ed77
          60792 => x"00", -- $0ed78
          60793 => x"00", -- $0ed79
          60794 => x"00", -- $0ed7a
          60795 => x"00", -- $0ed7b
          60796 => x"00", -- $0ed7c
          60797 => x"00", -- $0ed7d
          60798 => x"00", -- $0ed7e
          60799 => x"00", -- $0ed7f
          60800 => x"00", -- $0ed80
          60801 => x"00", -- $0ed81
          60802 => x"00", -- $0ed82
          60803 => x"00", -- $0ed83
          60804 => x"00", -- $0ed84
          60805 => x"00", -- $0ed85
          60806 => x"00", -- $0ed86
          60807 => x"00", -- $0ed87
          60808 => x"00", -- $0ed88
          60809 => x"00", -- $0ed89
          60810 => x"00", -- $0ed8a
          60811 => x"00", -- $0ed8b
          60812 => x"00", -- $0ed8c
          60813 => x"00", -- $0ed8d
          60814 => x"00", -- $0ed8e
          60815 => x"00", -- $0ed8f
          60816 => x"00", -- $0ed90
          60817 => x"00", -- $0ed91
          60818 => x"00", -- $0ed92
          60819 => x"00", -- $0ed93
          60820 => x"00", -- $0ed94
          60821 => x"00", -- $0ed95
          60822 => x"00", -- $0ed96
          60823 => x"00", -- $0ed97
          60824 => x"00", -- $0ed98
          60825 => x"00", -- $0ed99
          60826 => x"00", -- $0ed9a
          60827 => x"00", -- $0ed9b
          60828 => x"00", -- $0ed9c
          60829 => x"00", -- $0ed9d
          60830 => x"00", -- $0ed9e
          60831 => x"00", -- $0ed9f
          60832 => x"00", -- $0eda0
          60833 => x"00", -- $0eda1
          60834 => x"00", -- $0eda2
          60835 => x"00", -- $0eda3
          60836 => x"00", -- $0eda4
          60837 => x"00", -- $0eda5
          60838 => x"00", -- $0eda6
          60839 => x"00", -- $0eda7
          60840 => x"00", -- $0eda8
          60841 => x"00", -- $0eda9
          60842 => x"00", -- $0edaa
          60843 => x"00", -- $0edab
          60844 => x"00", -- $0edac
          60845 => x"00", -- $0edad
          60846 => x"00", -- $0edae
          60847 => x"00", -- $0edaf
          60848 => x"00", -- $0edb0
          60849 => x"00", -- $0edb1
          60850 => x"00", -- $0edb2
          60851 => x"00", -- $0edb3
          60852 => x"00", -- $0edb4
          60853 => x"00", -- $0edb5
          60854 => x"00", -- $0edb6
          60855 => x"00", -- $0edb7
          60856 => x"00", -- $0edb8
          60857 => x"00", -- $0edb9
          60858 => x"00", -- $0edba
          60859 => x"00", -- $0edbb
          60860 => x"00", -- $0edbc
          60861 => x"00", -- $0edbd
          60862 => x"00", -- $0edbe
          60863 => x"00", -- $0edbf
          60864 => x"00", -- $0edc0
          60865 => x"00", -- $0edc1
          60866 => x"00", -- $0edc2
          60867 => x"00", -- $0edc3
          60868 => x"00", -- $0edc4
          60869 => x"00", -- $0edc5
          60870 => x"00", -- $0edc6
          60871 => x"00", -- $0edc7
          60872 => x"00", -- $0edc8
          60873 => x"00", -- $0edc9
          60874 => x"00", -- $0edca
          60875 => x"00", -- $0edcb
          60876 => x"00", -- $0edcc
          60877 => x"00", -- $0edcd
          60878 => x"00", -- $0edce
          60879 => x"00", -- $0edcf
          60880 => x"00", -- $0edd0
          60881 => x"00", -- $0edd1
          60882 => x"00", -- $0edd2
          60883 => x"00", -- $0edd3
          60884 => x"00", -- $0edd4
          60885 => x"00", -- $0edd5
          60886 => x"00", -- $0edd6
          60887 => x"00", -- $0edd7
          60888 => x"00", -- $0edd8
          60889 => x"00", -- $0edd9
          60890 => x"00", -- $0edda
          60891 => x"00", -- $0eddb
          60892 => x"00", -- $0eddc
          60893 => x"00", -- $0eddd
          60894 => x"00", -- $0edde
          60895 => x"00", -- $0eddf
          60896 => x"00", -- $0ede0
          60897 => x"00", -- $0ede1
          60898 => x"00", -- $0ede2
          60899 => x"00", -- $0ede3
          60900 => x"00", -- $0ede4
          60901 => x"00", -- $0ede5
          60902 => x"00", -- $0ede6
          60903 => x"00", -- $0ede7
          60904 => x"00", -- $0ede8
          60905 => x"00", -- $0ede9
          60906 => x"00", -- $0edea
          60907 => x"00", -- $0edeb
          60908 => x"00", -- $0edec
          60909 => x"00", -- $0eded
          60910 => x"00", -- $0edee
          60911 => x"00", -- $0edef
          60912 => x"00", -- $0edf0
          60913 => x"00", -- $0edf1
          60914 => x"00", -- $0edf2
          60915 => x"00", -- $0edf3
          60916 => x"00", -- $0edf4
          60917 => x"00", -- $0edf5
          60918 => x"00", -- $0edf6
          60919 => x"00", -- $0edf7
          60920 => x"00", -- $0edf8
          60921 => x"00", -- $0edf9
          60922 => x"00", -- $0edfa
          60923 => x"00", -- $0edfb
          60924 => x"00", -- $0edfc
          60925 => x"00", -- $0edfd
          60926 => x"00", -- $0edfe
          60927 => x"00", -- $0edff
          60928 => x"00", -- $0ee00
          60929 => x"00", -- $0ee01
          60930 => x"00", -- $0ee02
          60931 => x"00", -- $0ee03
          60932 => x"00", -- $0ee04
          60933 => x"00", -- $0ee05
          60934 => x"00", -- $0ee06
          60935 => x"00", -- $0ee07
          60936 => x"00", -- $0ee08
          60937 => x"00", -- $0ee09
          60938 => x"00", -- $0ee0a
          60939 => x"00", -- $0ee0b
          60940 => x"00", -- $0ee0c
          60941 => x"00", -- $0ee0d
          60942 => x"00", -- $0ee0e
          60943 => x"00", -- $0ee0f
          60944 => x"00", -- $0ee10
          60945 => x"00", -- $0ee11
          60946 => x"00", -- $0ee12
          60947 => x"00", -- $0ee13
          60948 => x"00", -- $0ee14
          60949 => x"00", -- $0ee15
          60950 => x"00", -- $0ee16
          60951 => x"00", -- $0ee17
          60952 => x"00", -- $0ee18
          60953 => x"00", -- $0ee19
          60954 => x"00", -- $0ee1a
          60955 => x"00", -- $0ee1b
          60956 => x"00", -- $0ee1c
          60957 => x"00", -- $0ee1d
          60958 => x"00", -- $0ee1e
          60959 => x"00", -- $0ee1f
          60960 => x"00", -- $0ee20
          60961 => x"00", -- $0ee21
          60962 => x"00", -- $0ee22
          60963 => x"00", -- $0ee23
          60964 => x"00", -- $0ee24
          60965 => x"00", -- $0ee25
          60966 => x"00", -- $0ee26
          60967 => x"00", -- $0ee27
          60968 => x"00", -- $0ee28
          60969 => x"00", -- $0ee29
          60970 => x"00", -- $0ee2a
          60971 => x"00", -- $0ee2b
          60972 => x"00", -- $0ee2c
          60973 => x"00", -- $0ee2d
          60974 => x"00", -- $0ee2e
          60975 => x"00", -- $0ee2f
          60976 => x"00", -- $0ee30
          60977 => x"00", -- $0ee31
          60978 => x"00", -- $0ee32
          60979 => x"00", -- $0ee33
          60980 => x"00", -- $0ee34
          60981 => x"00", -- $0ee35
          60982 => x"00", -- $0ee36
          60983 => x"00", -- $0ee37
          60984 => x"00", -- $0ee38
          60985 => x"00", -- $0ee39
          60986 => x"00", -- $0ee3a
          60987 => x"00", -- $0ee3b
          60988 => x"00", -- $0ee3c
          60989 => x"00", -- $0ee3d
          60990 => x"00", -- $0ee3e
          60991 => x"00", -- $0ee3f
          60992 => x"00", -- $0ee40
          60993 => x"00", -- $0ee41
          60994 => x"00", -- $0ee42
          60995 => x"00", -- $0ee43
          60996 => x"00", -- $0ee44
          60997 => x"00", -- $0ee45
          60998 => x"00", -- $0ee46
          60999 => x"00", -- $0ee47
          61000 => x"00", -- $0ee48
          61001 => x"00", -- $0ee49
          61002 => x"00", -- $0ee4a
          61003 => x"00", -- $0ee4b
          61004 => x"00", -- $0ee4c
          61005 => x"00", -- $0ee4d
          61006 => x"00", -- $0ee4e
          61007 => x"00", -- $0ee4f
          61008 => x"00", -- $0ee50
          61009 => x"00", -- $0ee51
          61010 => x"00", -- $0ee52
          61011 => x"00", -- $0ee53
          61012 => x"00", -- $0ee54
          61013 => x"00", -- $0ee55
          61014 => x"00", -- $0ee56
          61015 => x"00", -- $0ee57
          61016 => x"00", -- $0ee58
          61017 => x"00", -- $0ee59
          61018 => x"00", -- $0ee5a
          61019 => x"00", -- $0ee5b
          61020 => x"00", -- $0ee5c
          61021 => x"00", -- $0ee5d
          61022 => x"00", -- $0ee5e
          61023 => x"00", -- $0ee5f
          61024 => x"00", -- $0ee60
          61025 => x"00", -- $0ee61
          61026 => x"00", -- $0ee62
          61027 => x"00", -- $0ee63
          61028 => x"00", -- $0ee64
          61029 => x"00", -- $0ee65
          61030 => x"00", -- $0ee66
          61031 => x"00", -- $0ee67
          61032 => x"00", -- $0ee68
          61033 => x"00", -- $0ee69
          61034 => x"00", -- $0ee6a
          61035 => x"00", -- $0ee6b
          61036 => x"00", -- $0ee6c
          61037 => x"00", -- $0ee6d
          61038 => x"00", -- $0ee6e
          61039 => x"00", -- $0ee6f
          61040 => x"00", -- $0ee70
          61041 => x"00", -- $0ee71
          61042 => x"00", -- $0ee72
          61043 => x"00", -- $0ee73
          61044 => x"00", -- $0ee74
          61045 => x"00", -- $0ee75
          61046 => x"00", -- $0ee76
          61047 => x"00", -- $0ee77
          61048 => x"00", -- $0ee78
          61049 => x"00", -- $0ee79
          61050 => x"00", -- $0ee7a
          61051 => x"00", -- $0ee7b
          61052 => x"00", -- $0ee7c
          61053 => x"00", -- $0ee7d
          61054 => x"00", -- $0ee7e
          61055 => x"00", -- $0ee7f
          61056 => x"00", -- $0ee80
          61057 => x"00", -- $0ee81
          61058 => x"00", -- $0ee82
          61059 => x"00", -- $0ee83
          61060 => x"00", -- $0ee84
          61061 => x"00", -- $0ee85
          61062 => x"00", -- $0ee86
          61063 => x"00", -- $0ee87
          61064 => x"00", -- $0ee88
          61065 => x"00", -- $0ee89
          61066 => x"00", -- $0ee8a
          61067 => x"00", -- $0ee8b
          61068 => x"00", -- $0ee8c
          61069 => x"00", -- $0ee8d
          61070 => x"00", -- $0ee8e
          61071 => x"00", -- $0ee8f
          61072 => x"00", -- $0ee90
          61073 => x"00", -- $0ee91
          61074 => x"00", -- $0ee92
          61075 => x"00", -- $0ee93
          61076 => x"00", -- $0ee94
          61077 => x"00", -- $0ee95
          61078 => x"00", -- $0ee96
          61079 => x"00", -- $0ee97
          61080 => x"00", -- $0ee98
          61081 => x"00", -- $0ee99
          61082 => x"00", -- $0ee9a
          61083 => x"00", -- $0ee9b
          61084 => x"00", -- $0ee9c
          61085 => x"00", -- $0ee9d
          61086 => x"00", -- $0ee9e
          61087 => x"00", -- $0ee9f
          61088 => x"00", -- $0eea0
          61089 => x"00", -- $0eea1
          61090 => x"00", -- $0eea2
          61091 => x"00", -- $0eea3
          61092 => x"00", -- $0eea4
          61093 => x"00", -- $0eea5
          61094 => x"00", -- $0eea6
          61095 => x"00", -- $0eea7
          61096 => x"00", -- $0eea8
          61097 => x"00", -- $0eea9
          61098 => x"00", -- $0eeaa
          61099 => x"00", -- $0eeab
          61100 => x"00", -- $0eeac
          61101 => x"00", -- $0eead
          61102 => x"00", -- $0eeae
          61103 => x"00", -- $0eeaf
          61104 => x"00", -- $0eeb0
          61105 => x"00", -- $0eeb1
          61106 => x"00", -- $0eeb2
          61107 => x"00", -- $0eeb3
          61108 => x"00", -- $0eeb4
          61109 => x"00", -- $0eeb5
          61110 => x"00", -- $0eeb6
          61111 => x"00", -- $0eeb7
          61112 => x"00", -- $0eeb8
          61113 => x"00", -- $0eeb9
          61114 => x"00", -- $0eeba
          61115 => x"00", -- $0eebb
          61116 => x"00", -- $0eebc
          61117 => x"00", -- $0eebd
          61118 => x"00", -- $0eebe
          61119 => x"00", -- $0eebf
          61120 => x"00", -- $0eec0
          61121 => x"00", -- $0eec1
          61122 => x"00", -- $0eec2
          61123 => x"00", -- $0eec3
          61124 => x"00", -- $0eec4
          61125 => x"00", -- $0eec5
          61126 => x"00", -- $0eec6
          61127 => x"00", -- $0eec7
          61128 => x"00", -- $0eec8
          61129 => x"00", -- $0eec9
          61130 => x"00", -- $0eeca
          61131 => x"00", -- $0eecb
          61132 => x"00", -- $0eecc
          61133 => x"00", -- $0eecd
          61134 => x"00", -- $0eece
          61135 => x"00", -- $0eecf
          61136 => x"00", -- $0eed0
          61137 => x"00", -- $0eed1
          61138 => x"00", -- $0eed2
          61139 => x"00", -- $0eed3
          61140 => x"00", -- $0eed4
          61141 => x"00", -- $0eed5
          61142 => x"00", -- $0eed6
          61143 => x"00", -- $0eed7
          61144 => x"00", -- $0eed8
          61145 => x"00", -- $0eed9
          61146 => x"00", -- $0eeda
          61147 => x"00", -- $0eedb
          61148 => x"00", -- $0eedc
          61149 => x"00", -- $0eedd
          61150 => x"00", -- $0eede
          61151 => x"00", -- $0eedf
          61152 => x"00", -- $0eee0
          61153 => x"00", -- $0eee1
          61154 => x"00", -- $0eee2
          61155 => x"00", -- $0eee3
          61156 => x"00", -- $0eee4
          61157 => x"00", -- $0eee5
          61158 => x"00", -- $0eee6
          61159 => x"00", -- $0eee7
          61160 => x"00", -- $0eee8
          61161 => x"00", -- $0eee9
          61162 => x"00", -- $0eeea
          61163 => x"00", -- $0eeeb
          61164 => x"00", -- $0eeec
          61165 => x"00", -- $0eeed
          61166 => x"00", -- $0eeee
          61167 => x"00", -- $0eeef
          61168 => x"00", -- $0eef0
          61169 => x"00", -- $0eef1
          61170 => x"00", -- $0eef2
          61171 => x"00", -- $0eef3
          61172 => x"00", -- $0eef4
          61173 => x"00", -- $0eef5
          61174 => x"00", -- $0eef6
          61175 => x"00", -- $0eef7
          61176 => x"00", -- $0eef8
          61177 => x"00", -- $0eef9
          61178 => x"00", -- $0eefa
          61179 => x"00", -- $0eefb
          61180 => x"00", -- $0eefc
          61181 => x"00", -- $0eefd
          61182 => x"00", -- $0eefe
          61183 => x"00", -- $0eeff
          61184 => x"00", -- $0ef00
          61185 => x"00", -- $0ef01
          61186 => x"00", -- $0ef02
          61187 => x"00", -- $0ef03
          61188 => x"00", -- $0ef04
          61189 => x"00", -- $0ef05
          61190 => x"00", -- $0ef06
          61191 => x"00", -- $0ef07
          61192 => x"00", -- $0ef08
          61193 => x"00", -- $0ef09
          61194 => x"00", -- $0ef0a
          61195 => x"00", -- $0ef0b
          61196 => x"00", -- $0ef0c
          61197 => x"00", -- $0ef0d
          61198 => x"00", -- $0ef0e
          61199 => x"00", -- $0ef0f
          61200 => x"00", -- $0ef10
          61201 => x"00", -- $0ef11
          61202 => x"00", -- $0ef12
          61203 => x"00", -- $0ef13
          61204 => x"00", -- $0ef14
          61205 => x"00", -- $0ef15
          61206 => x"00", -- $0ef16
          61207 => x"00", -- $0ef17
          61208 => x"00", -- $0ef18
          61209 => x"00", -- $0ef19
          61210 => x"00", -- $0ef1a
          61211 => x"00", -- $0ef1b
          61212 => x"00", -- $0ef1c
          61213 => x"00", -- $0ef1d
          61214 => x"00", -- $0ef1e
          61215 => x"00", -- $0ef1f
          61216 => x"00", -- $0ef20
          61217 => x"00", -- $0ef21
          61218 => x"00", -- $0ef22
          61219 => x"00", -- $0ef23
          61220 => x"00", -- $0ef24
          61221 => x"00", -- $0ef25
          61222 => x"00", -- $0ef26
          61223 => x"00", -- $0ef27
          61224 => x"00", -- $0ef28
          61225 => x"00", -- $0ef29
          61226 => x"00", -- $0ef2a
          61227 => x"00", -- $0ef2b
          61228 => x"00", -- $0ef2c
          61229 => x"00", -- $0ef2d
          61230 => x"00", -- $0ef2e
          61231 => x"00", -- $0ef2f
          61232 => x"00", -- $0ef30
          61233 => x"00", -- $0ef31
          61234 => x"00", -- $0ef32
          61235 => x"00", -- $0ef33
          61236 => x"00", -- $0ef34
          61237 => x"00", -- $0ef35
          61238 => x"00", -- $0ef36
          61239 => x"00", -- $0ef37
          61240 => x"00", -- $0ef38
          61241 => x"00", -- $0ef39
          61242 => x"00", -- $0ef3a
          61243 => x"00", -- $0ef3b
          61244 => x"00", -- $0ef3c
          61245 => x"00", -- $0ef3d
          61246 => x"00", -- $0ef3e
          61247 => x"00", -- $0ef3f
          61248 => x"00", -- $0ef40
          61249 => x"00", -- $0ef41
          61250 => x"00", -- $0ef42
          61251 => x"00", -- $0ef43
          61252 => x"00", -- $0ef44
          61253 => x"00", -- $0ef45
          61254 => x"00", -- $0ef46
          61255 => x"00", -- $0ef47
          61256 => x"00", -- $0ef48
          61257 => x"00", -- $0ef49
          61258 => x"00", -- $0ef4a
          61259 => x"00", -- $0ef4b
          61260 => x"00", -- $0ef4c
          61261 => x"00", -- $0ef4d
          61262 => x"00", -- $0ef4e
          61263 => x"00", -- $0ef4f
          61264 => x"00", -- $0ef50
          61265 => x"00", -- $0ef51
          61266 => x"00", -- $0ef52
          61267 => x"00", -- $0ef53
          61268 => x"00", -- $0ef54
          61269 => x"00", -- $0ef55
          61270 => x"00", -- $0ef56
          61271 => x"00", -- $0ef57
          61272 => x"00", -- $0ef58
          61273 => x"00", -- $0ef59
          61274 => x"00", -- $0ef5a
          61275 => x"00", -- $0ef5b
          61276 => x"00", -- $0ef5c
          61277 => x"00", -- $0ef5d
          61278 => x"00", -- $0ef5e
          61279 => x"00", -- $0ef5f
          61280 => x"00", -- $0ef60
          61281 => x"00", -- $0ef61
          61282 => x"00", -- $0ef62
          61283 => x"00", -- $0ef63
          61284 => x"00", -- $0ef64
          61285 => x"00", -- $0ef65
          61286 => x"00", -- $0ef66
          61287 => x"00", -- $0ef67
          61288 => x"00", -- $0ef68
          61289 => x"00", -- $0ef69
          61290 => x"00", -- $0ef6a
          61291 => x"00", -- $0ef6b
          61292 => x"00", -- $0ef6c
          61293 => x"00", -- $0ef6d
          61294 => x"00", -- $0ef6e
          61295 => x"00", -- $0ef6f
          61296 => x"00", -- $0ef70
          61297 => x"00", -- $0ef71
          61298 => x"00", -- $0ef72
          61299 => x"00", -- $0ef73
          61300 => x"00", -- $0ef74
          61301 => x"00", -- $0ef75
          61302 => x"00", -- $0ef76
          61303 => x"00", -- $0ef77
          61304 => x"00", -- $0ef78
          61305 => x"00", -- $0ef79
          61306 => x"00", -- $0ef7a
          61307 => x"00", -- $0ef7b
          61308 => x"00", -- $0ef7c
          61309 => x"00", -- $0ef7d
          61310 => x"00", -- $0ef7e
          61311 => x"00", -- $0ef7f
          61312 => x"00", -- $0ef80
          61313 => x"00", -- $0ef81
          61314 => x"00", -- $0ef82
          61315 => x"00", -- $0ef83
          61316 => x"00", -- $0ef84
          61317 => x"00", -- $0ef85
          61318 => x"00", -- $0ef86
          61319 => x"00", -- $0ef87
          61320 => x"00", -- $0ef88
          61321 => x"00", -- $0ef89
          61322 => x"00", -- $0ef8a
          61323 => x"00", -- $0ef8b
          61324 => x"00", -- $0ef8c
          61325 => x"00", -- $0ef8d
          61326 => x"00", -- $0ef8e
          61327 => x"00", -- $0ef8f
          61328 => x"00", -- $0ef90
          61329 => x"00", -- $0ef91
          61330 => x"00", -- $0ef92
          61331 => x"00", -- $0ef93
          61332 => x"00", -- $0ef94
          61333 => x"00", -- $0ef95
          61334 => x"00", -- $0ef96
          61335 => x"00", -- $0ef97
          61336 => x"00", -- $0ef98
          61337 => x"00", -- $0ef99
          61338 => x"00", -- $0ef9a
          61339 => x"00", -- $0ef9b
          61340 => x"00", -- $0ef9c
          61341 => x"00", -- $0ef9d
          61342 => x"00", -- $0ef9e
          61343 => x"00", -- $0ef9f
          61344 => x"00", -- $0efa0
          61345 => x"00", -- $0efa1
          61346 => x"00", -- $0efa2
          61347 => x"00", -- $0efa3
          61348 => x"00", -- $0efa4
          61349 => x"00", -- $0efa5
          61350 => x"00", -- $0efa6
          61351 => x"00", -- $0efa7
          61352 => x"00", -- $0efa8
          61353 => x"00", -- $0efa9
          61354 => x"00", -- $0efaa
          61355 => x"00", -- $0efab
          61356 => x"00", -- $0efac
          61357 => x"00", -- $0efad
          61358 => x"00", -- $0efae
          61359 => x"00", -- $0efaf
          61360 => x"00", -- $0efb0
          61361 => x"00", -- $0efb1
          61362 => x"00", -- $0efb2
          61363 => x"00", -- $0efb3
          61364 => x"00", -- $0efb4
          61365 => x"00", -- $0efb5
          61366 => x"00", -- $0efb6
          61367 => x"00", -- $0efb7
          61368 => x"00", -- $0efb8
          61369 => x"00", -- $0efb9
          61370 => x"00", -- $0efba
          61371 => x"00", -- $0efbb
          61372 => x"00", -- $0efbc
          61373 => x"00", -- $0efbd
          61374 => x"00", -- $0efbe
          61375 => x"00", -- $0efbf
          61376 => x"00", -- $0efc0
          61377 => x"00", -- $0efc1
          61378 => x"00", -- $0efc2
          61379 => x"00", -- $0efc3
          61380 => x"00", -- $0efc4
          61381 => x"00", -- $0efc5
          61382 => x"00", -- $0efc6
          61383 => x"00", -- $0efc7
          61384 => x"00", -- $0efc8
          61385 => x"00", -- $0efc9
          61386 => x"00", -- $0efca
          61387 => x"00", -- $0efcb
          61388 => x"00", -- $0efcc
          61389 => x"00", -- $0efcd
          61390 => x"00", -- $0efce
          61391 => x"00", -- $0efcf
          61392 => x"00", -- $0efd0
          61393 => x"00", -- $0efd1
          61394 => x"00", -- $0efd2
          61395 => x"00", -- $0efd3
          61396 => x"00", -- $0efd4
          61397 => x"00", -- $0efd5
          61398 => x"00", -- $0efd6
          61399 => x"00", -- $0efd7
          61400 => x"00", -- $0efd8
          61401 => x"00", -- $0efd9
          61402 => x"00", -- $0efda
          61403 => x"00", -- $0efdb
          61404 => x"00", -- $0efdc
          61405 => x"00", -- $0efdd
          61406 => x"00", -- $0efde
          61407 => x"00", -- $0efdf
          61408 => x"00", -- $0efe0
          61409 => x"00", -- $0efe1
          61410 => x"00", -- $0efe2
          61411 => x"00", -- $0efe3
          61412 => x"00", -- $0efe4
          61413 => x"00", -- $0efe5
          61414 => x"00", -- $0efe6
          61415 => x"00", -- $0efe7
          61416 => x"00", -- $0efe8
          61417 => x"00", -- $0efe9
          61418 => x"00", -- $0efea
          61419 => x"00", -- $0efeb
          61420 => x"00", -- $0efec
          61421 => x"00", -- $0efed
          61422 => x"00", -- $0efee
          61423 => x"00", -- $0efef
          61424 => x"00", -- $0eff0
          61425 => x"00", -- $0eff1
          61426 => x"00", -- $0eff2
          61427 => x"00", -- $0eff3
          61428 => x"00", -- $0eff4
          61429 => x"00", -- $0eff5
          61430 => x"00", -- $0eff6
          61431 => x"00", -- $0eff7
          61432 => x"00", -- $0eff8
          61433 => x"00", -- $0eff9
          61434 => x"00", -- $0effa
          61435 => x"00", -- $0effb
          61436 => x"00", -- $0effc
          61437 => x"00", -- $0effd
          61438 => x"00", -- $0effe
          61439 => x"00", -- $0efff
          61440 => x"00", -- $0f000
          61441 => x"00", -- $0f001
          61442 => x"00", -- $0f002
          61443 => x"00", -- $0f003
          61444 => x"00", -- $0f004
          61445 => x"00", -- $0f005
          61446 => x"00", -- $0f006
          61447 => x"00", -- $0f007
          61448 => x"00", -- $0f008
          61449 => x"00", -- $0f009
          61450 => x"00", -- $0f00a
          61451 => x"00", -- $0f00b
          61452 => x"00", -- $0f00c
          61453 => x"00", -- $0f00d
          61454 => x"00", -- $0f00e
          61455 => x"00", -- $0f00f
          61456 => x"00", -- $0f010
          61457 => x"00", -- $0f011
          61458 => x"00", -- $0f012
          61459 => x"00", -- $0f013
          61460 => x"00", -- $0f014
          61461 => x"00", -- $0f015
          61462 => x"00", -- $0f016
          61463 => x"00", -- $0f017
          61464 => x"00", -- $0f018
          61465 => x"00", -- $0f019
          61466 => x"00", -- $0f01a
          61467 => x"00", -- $0f01b
          61468 => x"00", -- $0f01c
          61469 => x"00", -- $0f01d
          61470 => x"00", -- $0f01e
          61471 => x"00", -- $0f01f
          61472 => x"00", -- $0f020
          61473 => x"00", -- $0f021
          61474 => x"00", -- $0f022
          61475 => x"00", -- $0f023
          61476 => x"00", -- $0f024
          61477 => x"00", -- $0f025
          61478 => x"00", -- $0f026
          61479 => x"00", -- $0f027
          61480 => x"00", -- $0f028
          61481 => x"00", -- $0f029
          61482 => x"00", -- $0f02a
          61483 => x"00", -- $0f02b
          61484 => x"00", -- $0f02c
          61485 => x"00", -- $0f02d
          61486 => x"00", -- $0f02e
          61487 => x"00", -- $0f02f
          61488 => x"00", -- $0f030
          61489 => x"00", -- $0f031
          61490 => x"00", -- $0f032
          61491 => x"00", -- $0f033
          61492 => x"00", -- $0f034
          61493 => x"00", -- $0f035
          61494 => x"00", -- $0f036
          61495 => x"00", -- $0f037
          61496 => x"00", -- $0f038
          61497 => x"00", -- $0f039
          61498 => x"00", -- $0f03a
          61499 => x"00", -- $0f03b
          61500 => x"00", -- $0f03c
          61501 => x"00", -- $0f03d
          61502 => x"00", -- $0f03e
          61503 => x"00", -- $0f03f
          61504 => x"00", -- $0f040
          61505 => x"00", -- $0f041
          61506 => x"00", -- $0f042
          61507 => x"00", -- $0f043
          61508 => x"00", -- $0f044
          61509 => x"00", -- $0f045
          61510 => x"00", -- $0f046
          61511 => x"00", -- $0f047
          61512 => x"00", -- $0f048
          61513 => x"00", -- $0f049
          61514 => x"00", -- $0f04a
          61515 => x"00", -- $0f04b
          61516 => x"00", -- $0f04c
          61517 => x"00", -- $0f04d
          61518 => x"00", -- $0f04e
          61519 => x"00", -- $0f04f
          61520 => x"00", -- $0f050
          61521 => x"00", -- $0f051
          61522 => x"00", -- $0f052
          61523 => x"00", -- $0f053
          61524 => x"00", -- $0f054
          61525 => x"00", -- $0f055
          61526 => x"00", -- $0f056
          61527 => x"00", -- $0f057
          61528 => x"00", -- $0f058
          61529 => x"00", -- $0f059
          61530 => x"00", -- $0f05a
          61531 => x"00", -- $0f05b
          61532 => x"00", -- $0f05c
          61533 => x"00", -- $0f05d
          61534 => x"00", -- $0f05e
          61535 => x"00", -- $0f05f
          61536 => x"00", -- $0f060
          61537 => x"00", -- $0f061
          61538 => x"00", -- $0f062
          61539 => x"00", -- $0f063
          61540 => x"00", -- $0f064
          61541 => x"00", -- $0f065
          61542 => x"00", -- $0f066
          61543 => x"00", -- $0f067
          61544 => x"00", -- $0f068
          61545 => x"00", -- $0f069
          61546 => x"00", -- $0f06a
          61547 => x"00", -- $0f06b
          61548 => x"00", -- $0f06c
          61549 => x"00", -- $0f06d
          61550 => x"00", -- $0f06e
          61551 => x"00", -- $0f06f
          61552 => x"00", -- $0f070
          61553 => x"00", -- $0f071
          61554 => x"00", -- $0f072
          61555 => x"00", -- $0f073
          61556 => x"00", -- $0f074
          61557 => x"00", -- $0f075
          61558 => x"00", -- $0f076
          61559 => x"00", -- $0f077
          61560 => x"00", -- $0f078
          61561 => x"00", -- $0f079
          61562 => x"00", -- $0f07a
          61563 => x"00", -- $0f07b
          61564 => x"00", -- $0f07c
          61565 => x"00", -- $0f07d
          61566 => x"00", -- $0f07e
          61567 => x"00", -- $0f07f
          61568 => x"00", -- $0f080
          61569 => x"00", -- $0f081
          61570 => x"00", -- $0f082
          61571 => x"00", -- $0f083
          61572 => x"00", -- $0f084
          61573 => x"00", -- $0f085
          61574 => x"00", -- $0f086
          61575 => x"00", -- $0f087
          61576 => x"00", -- $0f088
          61577 => x"00", -- $0f089
          61578 => x"00", -- $0f08a
          61579 => x"00", -- $0f08b
          61580 => x"00", -- $0f08c
          61581 => x"00", -- $0f08d
          61582 => x"00", -- $0f08e
          61583 => x"00", -- $0f08f
          61584 => x"00", -- $0f090
          61585 => x"00", -- $0f091
          61586 => x"00", -- $0f092
          61587 => x"00", -- $0f093
          61588 => x"00", -- $0f094
          61589 => x"00", -- $0f095
          61590 => x"00", -- $0f096
          61591 => x"00", -- $0f097
          61592 => x"00", -- $0f098
          61593 => x"00", -- $0f099
          61594 => x"00", -- $0f09a
          61595 => x"00", -- $0f09b
          61596 => x"00", -- $0f09c
          61597 => x"00", -- $0f09d
          61598 => x"00", -- $0f09e
          61599 => x"00", -- $0f09f
          61600 => x"00", -- $0f0a0
          61601 => x"00", -- $0f0a1
          61602 => x"00", -- $0f0a2
          61603 => x"00", -- $0f0a3
          61604 => x"00", -- $0f0a4
          61605 => x"00", -- $0f0a5
          61606 => x"00", -- $0f0a6
          61607 => x"00", -- $0f0a7
          61608 => x"00", -- $0f0a8
          61609 => x"00", -- $0f0a9
          61610 => x"00", -- $0f0aa
          61611 => x"00", -- $0f0ab
          61612 => x"00", -- $0f0ac
          61613 => x"00", -- $0f0ad
          61614 => x"00", -- $0f0ae
          61615 => x"00", -- $0f0af
          61616 => x"00", -- $0f0b0
          61617 => x"00", -- $0f0b1
          61618 => x"00", -- $0f0b2
          61619 => x"00", -- $0f0b3
          61620 => x"00", -- $0f0b4
          61621 => x"00", -- $0f0b5
          61622 => x"00", -- $0f0b6
          61623 => x"00", -- $0f0b7
          61624 => x"00", -- $0f0b8
          61625 => x"00", -- $0f0b9
          61626 => x"00", -- $0f0ba
          61627 => x"00", -- $0f0bb
          61628 => x"00", -- $0f0bc
          61629 => x"00", -- $0f0bd
          61630 => x"00", -- $0f0be
          61631 => x"00", -- $0f0bf
          61632 => x"00", -- $0f0c0
          61633 => x"00", -- $0f0c1
          61634 => x"00", -- $0f0c2
          61635 => x"00", -- $0f0c3
          61636 => x"00", -- $0f0c4
          61637 => x"00", -- $0f0c5
          61638 => x"00", -- $0f0c6
          61639 => x"00", -- $0f0c7
          61640 => x"00", -- $0f0c8
          61641 => x"00", -- $0f0c9
          61642 => x"00", -- $0f0ca
          61643 => x"00", -- $0f0cb
          61644 => x"00", -- $0f0cc
          61645 => x"00", -- $0f0cd
          61646 => x"00", -- $0f0ce
          61647 => x"00", -- $0f0cf
          61648 => x"00", -- $0f0d0
          61649 => x"00", -- $0f0d1
          61650 => x"00", -- $0f0d2
          61651 => x"00", -- $0f0d3
          61652 => x"00", -- $0f0d4
          61653 => x"00", -- $0f0d5
          61654 => x"00", -- $0f0d6
          61655 => x"00", -- $0f0d7
          61656 => x"00", -- $0f0d8
          61657 => x"00", -- $0f0d9
          61658 => x"00", -- $0f0da
          61659 => x"00", -- $0f0db
          61660 => x"00", -- $0f0dc
          61661 => x"00", -- $0f0dd
          61662 => x"00", -- $0f0de
          61663 => x"00", -- $0f0df
          61664 => x"00", -- $0f0e0
          61665 => x"00", -- $0f0e1
          61666 => x"00", -- $0f0e2
          61667 => x"00", -- $0f0e3
          61668 => x"00", -- $0f0e4
          61669 => x"00", -- $0f0e5
          61670 => x"00", -- $0f0e6
          61671 => x"00", -- $0f0e7
          61672 => x"00", -- $0f0e8
          61673 => x"00", -- $0f0e9
          61674 => x"00", -- $0f0ea
          61675 => x"00", -- $0f0eb
          61676 => x"00", -- $0f0ec
          61677 => x"00", -- $0f0ed
          61678 => x"00", -- $0f0ee
          61679 => x"00", -- $0f0ef
          61680 => x"00", -- $0f0f0
          61681 => x"00", -- $0f0f1
          61682 => x"00", -- $0f0f2
          61683 => x"00", -- $0f0f3
          61684 => x"00", -- $0f0f4
          61685 => x"00", -- $0f0f5
          61686 => x"00", -- $0f0f6
          61687 => x"00", -- $0f0f7
          61688 => x"00", -- $0f0f8
          61689 => x"00", -- $0f0f9
          61690 => x"00", -- $0f0fa
          61691 => x"00", -- $0f0fb
          61692 => x"00", -- $0f0fc
          61693 => x"00", -- $0f0fd
          61694 => x"00", -- $0f0fe
          61695 => x"00", -- $0f0ff
          61696 => x"00", -- $0f100
          61697 => x"00", -- $0f101
          61698 => x"00", -- $0f102
          61699 => x"00", -- $0f103
          61700 => x"00", -- $0f104
          61701 => x"00", -- $0f105
          61702 => x"00", -- $0f106
          61703 => x"00", -- $0f107
          61704 => x"00", -- $0f108
          61705 => x"00", -- $0f109
          61706 => x"00", -- $0f10a
          61707 => x"00", -- $0f10b
          61708 => x"00", -- $0f10c
          61709 => x"00", -- $0f10d
          61710 => x"00", -- $0f10e
          61711 => x"00", -- $0f10f
          61712 => x"00", -- $0f110
          61713 => x"00", -- $0f111
          61714 => x"00", -- $0f112
          61715 => x"00", -- $0f113
          61716 => x"00", -- $0f114
          61717 => x"00", -- $0f115
          61718 => x"00", -- $0f116
          61719 => x"00", -- $0f117
          61720 => x"00", -- $0f118
          61721 => x"00", -- $0f119
          61722 => x"00", -- $0f11a
          61723 => x"00", -- $0f11b
          61724 => x"00", -- $0f11c
          61725 => x"00", -- $0f11d
          61726 => x"00", -- $0f11e
          61727 => x"00", -- $0f11f
          61728 => x"00", -- $0f120
          61729 => x"00", -- $0f121
          61730 => x"00", -- $0f122
          61731 => x"00", -- $0f123
          61732 => x"00", -- $0f124
          61733 => x"00", -- $0f125
          61734 => x"00", -- $0f126
          61735 => x"00", -- $0f127
          61736 => x"00", -- $0f128
          61737 => x"00", -- $0f129
          61738 => x"00", -- $0f12a
          61739 => x"00", -- $0f12b
          61740 => x"00", -- $0f12c
          61741 => x"00", -- $0f12d
          61742 => x"00", -- $0f12e
          61743 => x"00", -- $0f12f
          61744 => x"00", -- $0f130
          61745 => x"00", -- $0f131
          61746 => x"00", -- $0f132
          61747 => x"00", -- $0f133
          61748 => x"00", -- $0f134
          61749 => x"00", -- $0f135
          61750 => x"00", -- $0f136
          61751 => x"00", -- $0f137
          61752 => x"00", -- $0f138
          61753 => x"00", -- $0f139
          61754 => x"00", -- $0f13a
          61755 => x"00", -- $0f13b
          61756 => x"00", -- $0f13c
          61757 => x"00", -- $0f13d
          61758 => x"00", -- $0f13e
          61759 => x"00", -- $0f13f
          61760 => x"00", -- $0f140
          61761 => x"00", -- $0f141
          61762 => x"00", -- $0f142
          61763 => x"00", -- $0f143
          61764 => x"00", -- $0f144
          61765 => x"00", -- $0f145
          61766 => x"00", -- $0f146
          61767 => x"00", -- $0f147
          61768 => x"00", -- $0f148
          61769 => x"00", -- $0f149
          61770 => x"00", -- $0f14a
          61771 => x"00", -- $0f14b
          61772 => x"00", -- $0f14c
          61773 => x"00", -- $0f14d
          61774 => x"00", -- $0f14e
          61775 => x"00", -- $0f14f
          61776 => x"00", -- $0f150
          61777 => x"00", -- $0f151
          61778 => x"00", -- $0f152
          61779 => x"00", -- $0f153
          61780 => x"00", -- $0f154
          61781 => x"00", -- $0f155
          61782 => x"00", -- $0f156
          61783 => x"00", -- $0f157
          61784 => x"00", -- $0f158
          61785 => x"00", -- $0f159
          61786 => x"00", -- $0f15a
          61787 => x"00", -- $0f15b
          61788 => x"00", -- $0f15c
          61789 => x"00", -- $0f15d
          61790 => x"00", -- $0f15e
          61791 => x"00", -- $0f15f
          61792 => x"00", -- $0f160
          61793 => x"00", -- $0f161
          61794 => x"00", -- $0f162
          61795 => x"00", -- $0f163
          61796 => x"00", -- $0f164
          61797 => x"00", -- $0f165
          61798 => x"00", -- $0f166
          61799 => x"00", -- $0f167
          61800 => x"00", -- $0f168
          61801 => x"00", -- $0f169
          61802 => x"00", -- $0f16a
          61803 => x"00", -- $0f16b
          61804 => x"00", -- $0f16c
          61805 => x"00", -- $0f16d
          61806 => x"00", -- $0f16e
          61807 => x"00", -- $0f16f
          61808 => x"00", -- $0f170
          61809 => x"00", -- $0f171
          61810 => x"00", -- $0f172
          61811 => x"00", -- $0f173
          61812 => x"00", -- $0f174
          61813 => x"00", -- $0f175
          61814 => x"00", -- $0f176
          61815 => x"00", -- $0f177
          61816 => x"00", -- $0f178
          61817 => x"00", -- $0f179
          61818 => x"00", -- $0f17a
          61819 => x"00", -- $0f17b
          61820 => x"00", -- $0f17c
          61821 => x"00", -- $0f17d
          61822 => x"00", -- $0f17e
          61823 => x"00", -- $0f17f
          61824 => x"00", -- $0f180
          61825 => x"00", -- $0f181
          61826 => x"00", -- $0f182
          61827 => x"00", -- $0f183
          61828 => x"00", -- $0f184
          61829 => x"00", -- $0f185
          61830 => x"00", -- $0f186
          61831 => x"00", -- $0f187
          61832 => x"00", -- $0f188
          61833 => x"00", -- $0f189
          61834 => x"00", -- $0f18a
          61835 => x"00", -- $0f18b
          61836 => x"00", -- $0f18c
          61837 => x"00", -- $0f18d
          61838 => x"00", -- $0f18e
          61839 => x"00", -- $0f18f
          61840 => x"00", -- $0f190
          61841 => x"00", -- $0f191
          61842 => x"00", -- $0f192
          61843 => x"00", -- $0f193
          61844 => x"00", -- $0f194
          61845 => x"00", -- $0f195
          61846 => x"00", -- $0f196
          61847 => x"00", -- $0f197
          61848 => x"00", -- $0f198
          61849 => x"00", -- $0f199
          61850 => x"00", -- $0f19a
          61851 => x"00", -- $0f19b
          61852 => x"00", -- $0f19c
          61853 => x"00", -- $0f19d
          61854 => x"00", -- $0f19e
          61855 => x"00", -- $0f19f
          61856 => x"00", -- $0f1a0
          61857 => x"00", -- $0f1a1
          61858 => x"00", -- $0f1a2
          61859 => x"00", -- $0f1a3
          61860 => x"00", -- $0f1a4
          61861 => x"00", -- $0f1a5
          61862 => x"00", -- $0f1a6
          61863 => x"00", -- $0f1a7
          61864 => x"00", -- $0f1a8
          61865 => x"00", -- $0f1a9
          61866 => x"00", -- $0f1aa
          61867 => x"00", -- $0f1ab
          61868 => x"00", -- $0f1ac
          61869 => x"00", -- $0f1ad
          61870 => x"00", -- $0f1ae
          61871 => x"00", -- $0f1af
          61872 => x"00", -- $0f1b0
          61873 => x"00", -- $0f1b1
          61874 => x"00", -- $0f1b2
          61875 => x"00", -- $0f1b3
          61876 => x"00", -- $0f1b4
          61877 => x"00", -- $0f1b5
          61878 => x"00", -- $0f1b6
          61879 => x"00", -- $0f1b7
          61880 => x"00", -- $0f1b8
          61881 => x"00", -- $0f1b9
          61882 => x"00", -- $0f1ba
          61883 => x"00", -- $0f1bb
          61884 => x"00", -- $0f1bc
          61885 => x"00", -- $0f1bd
          61886 => x"00", -- $0f1be
          61887 => x"00", -- $0f1bf
          61888 => x"00", -- $0f1c0
          61889 => x"00", -- $0f1c1
          61890 => x"00", -- $0f1c2
          61891 => x"00", -- $0f1c3
          61892 => x"00", -- $0f1c4
          61893 => x"00", -- $0f1c5
          61894 => x"00", -- $0f1c6
          61895 => x"00", -- $0f1c7
          61896 => x"00", -- $0f1c8
          61897 => x"00", -- $0f1c9
          61898 => x"00", -- $0f1ca
          61899 => x"00", -- $0f1cb
          61900 => x"00", -- $0f1cc
          61901 => x"00", -- $0f1cd
          61902 => x"00", -- $0f1ce
          61903 => x"00", -- $0f1cf
          61904 => x"00", -- $0f1d0
          61905 => x"00", -- $0f1d1
          61906 => x"00", -- $0f1d2
          61907 => x"00", -- $0f1d3
          61908 => x"00", -- $0f1d4
          61909 => x"00", -- $0f1d5
          61910 => x"00", -- $0f1d6
          61911 => x"00", -- $0f1d7
          61912 => x"00", -- $0f1d8
          61913 => x"00", -- $0f1d9
          61914 => x"00", -- $0f1da
          61915 => x"00", -- $0f1db
          61916 => x"00", -- $0f1dc
          61917 => x"00", -- $0f1dd
          61918 => x"00", -- $0f1de
          61919 => x"00", -- $0f1df
          61920 => x"00", -- $0f1e0
          61921 => x"00", -- $0f1e1
          61922 => x"00", -- $0f1e2
          61923 => x"00", -- $0f1e3
          61924 => x"00", -- $0f1e4
          61925 => x"00", -- $0f1e5
          61926 => x"00", -- $0f1e6
          61927 => x"00", -- $0f1e7
          61928 => x"00", -- $0f1e8
          61929 => x"00", -- $0f1e9
          61930 => x"00", -- $0f1ea
          61931 => x"00", -- $0f1eb
          61932 => x"00", -- $0f1ec
          61933 => x"00", -- $0f1ed
          61934 => x"00", -- $0f1ee
          61935 => x"00", -- $0f1ef
          61936 => x"00", -- $0f1f0
          61937 => x"00", -- $0f1f1
          61938 => x"00", -- $0f1f2
          61939 => x"00", -- $0f1f3
          61940 => x"00", -- $0f1f4
          61941 => x"00", -- $0f1f5
          61942 => x"00", -- $0f1f6
          61943 => x"00", -- $0f1f7
          61944 => x"00", -- $0f1f8
          61945 => x"00", -- $0f1f9
          61946 => x"00", -- $0f1fa
          61947 => x"00", -- $0f1fb
          61948 => x"00", -- $0f1fc
          61949 => x"00", -- $0f1fd
          61950 => x"00", -- $0f1fe
          61951 => x"00", -- $0f1ff
          61952 => x"00", -- $0f200
          61953 => x"00", -- $0f201
          61954 => x"00", -- $0f202
          61955 => x"00", -- $0f203
          61956 => x"00", -- $0f204
          61957 => x"00", -- $0f205
          61958 => x"00", -- $0f206
          61959 => x"00", -- $0f207
          61960 => x"00", -- $0f208
          61961 => x"00", -- $0f209
          61962 => x"00", -- $0f20a
          61963 => x"00", -- $0f20b
          61964 => x"00", -- $0f20c
          61965 => x"00", -- $0f20d
          61966 => x"00", -- $0f20e
          61967 => x"00", -- $0f20f
          61968 => x"00", -- $0f210
          61969 => x"00", -- $0f211
          61970 => x"00", -- $0f212
          61971 => x"00", -- $0f213
          61972 => x"00", -- $0f214
          61973 => x"00", -- $0f215
          61974 => x"00", -- $0f216
          61975 => x"00", -- $0f217
          61976 => x"00", -- $0f218
          61977 => x"00", -- $0f219
          61978 => x"00", -- $0f21a
          61979 => x"00", -- $0f21b
          61980 => x"00", -- $0f21c
          61981 => x"00", -- $0f21d
          61982 => x"00", -- $0f21e
          61983 => x"00", -- $0f21f
          61984 => x"00", -- $0f220
          61985 => x"00", -- $0f221
          61986 => x"00", -- $0f222
          61987 => x"00", -- $0f223
          61988 => x"00", -- $0f224
          61989 => x"00", -- $0f225
          61990 => x"00", -- $0f226
          61991 => x"00", -- $0f227
          61992 => x"00", -- $0f228
          61993 => x"00", -- $0f229
          61994 => x"00", -- $0f22a
          61995 => x"00", -- $0f22b
          61996 => x"00", -- $0f22c
          61997 => x"00", -- $0f22d
          61998 => x"00", -- $0f22e
          61999 => x"00", -- $0f22f
          62000 => x"00", -- $0f230
          62001 => x"00", -- $0f231
          62002 => x"00", -- $0f232
          62003 => x"00", -- $0f233
          62004 => x"00", -- $0f234
          62005 => x"00", -- $0f235
          62006 => x"00", -- $0f236
          62007 => x"00", -- $0f237
          62008 => x"00", -- $0f238
          62009 => x"00", -- $0f239
          62010 => x"00", -- $0f23a
          62011 => x"00", -- $0f23b
          62012 => x"00", -- $0f23c
          62013 => x"00", -- $0f23d
          62014 => x"00", -- $0f23e
          62015 => x"00", -- $0f23f
          62016 => x"00", -- $0f240
          62017 => x"00", -- $0f241
          62018 => x"00", -- $0f242
          62019 => x"00", -- $0f243
          62020 => x"00", -- $0f244
          62021 => x"00", -- $0f245
          62022 => x"00", -- $0f246
          62023 => x"00", -- $0f247
          62024 => x"00", -- $0f248
          62025 => x"00", -- $0f249
          62026 => x"00", -- $0f24a
          62027 => x"00", -- $0f24b
          62028 => x"00", -- $0f24c
          62029 => x"00", -- $0f24d
          62030 => x"00", -- $0f24e
          62031 => x"00", -- $0f24f
          62032 => x"00", -- $0f250
          62033 => x"00", -- $0f251
          62034 => x"00", -- $0f252
          62035 => x"00", -- $0f253
          62036 => x"00", -- $0f254
          62037 => x"00", -- $0f255
          62038 => x"00", -- $0f256
          62039 => x"00", -- $0f257
          62040 => x"00", -- $0f258
          62041 => x"00", -- $0f259
          62042 => x"00", -- $0f25a
          62043 => x"00", -- $0f25b
          62044 => x"00", -- $0f25c
          62045 => x"00", -- $0f25d
          62046 => x"00", -- $0f25e
          62047 => x"00", -- $0f25f
          62048 => x"00", -- $0f260
          62049 => x"00", -- $0f261
          62050 => x"00", -- $0f262
          62051 => x"00", -- $0f263
          62052 => x"00", -- $0f264
          62053 => x"00", -- $0f265
          62054 => x"00", -- $0f266
          62055 => x"00", -- $0f267
          62056 => x"00", -- $0f268
          62057 => x"00", -- $0f269
          62058 => x"00", -- $0f26a
          62059 => x"00", -- $0f26b
          62060 => x"00", -- $0f26c
          62061 => x"00", -- $0f26d
          62062 => x"00", -- $0f26e
          62063 => x"00", -- $0f26f
          62064 => x"00", -- $0f270
          62065 => x"00", -- $0f271
          62066 => x"00", -- $0f272
          62067 => x"00", -- $0f273
          62068 => x"00", -- $0f274
          62069 => x"00", -- $0f275
          62070 => x"00", -- $0f276
          62071 => x"00", -- $0f277
          62072 => x"00", -- $0f278
          62073 => x"00", -- $0f279
          62074 => x"00", -- $0f27a
          62075 => x"00", -- $0f27b
          62076 => x"00", -- $0f27c
          62077 => x"00", -- $0f27d
          62078 => x"00", -- $0f27e
          62079 => x"00", -- $0f27f
          62080 => x"00", -- $0f280
          62081 => x"00", -- $0f281
          62082 => x"00", -- $0f282
          62083 => x"00", -- $0f283
          62084 => x"00", -- $0f284
          62085 => x"00", -- $0f285
          62086 => x"00", -- $0f286
          62087 => x"00", -- $0f287
          62088 => x"00", -- $0f288
          62089 => x"00", -- $0f289
          62090 => x"00", -- $0f28a
          62091 => x"00", -- $0f28b
          62092 => x"00", -- $0f28c
          62093 => x"00", -- $0f28d
          62094 => x"00", -- $0f28e
          62095 => x"00", -- $0f28f
          62096 => x"00", -- $0f290
          62097 => x"00", -- $0f291
          62098 => x"00", -- $0f292
          62099 => x"00", -- $0f293
          62100 => x"00", -- $0f294
          62101 => x"00", -- $0f295
          62102 => x"00", -- $0f296
          62103 => x"00", -- $0f297
          62104 => x"00", -- $0f298
          62105 => x"00", -- $0f299
          62106 => x"00", -- $0f29a
          62107 => x"00", -- $0f29b
          62108 => x"00", -- $0f29c
          62109 => x"00", -- $0f29d
          62110 => x"00", -- $0f29e
          62111 => x"00", -- $0f29f
          62112 => x"00", -- $0f2a0
          62113 => x"00", -- $0f2a1
          62114 => x"00", -- $0f2a2
          62115 => x"00", -- $0f2a3
          62116 => x"00", -- $0f2a4
          62117 => x"00", -- $0f2a5
          62118 => x"00", -- $0f2a6
          62119 => x"00", -- $0f2a7
          62120 => x"00", -- $0f2a8
          62121 => x"00", -- $0f2a9
          62122 => x"00", -- $0f2aa
          62123 => x"00", -- $0f2ab
          62124 => x"00", -- $0f2ac
          62125 => x"00", -- $0f2ad
          62126 => x"00", -- $0f2ae
          62127 => x"00", -- $0f2af
          62128 => x"00", -- $0f2b0
          62129 => x"00", -- $0f2b1
          62130 => x"00", -- $0f2b2
          62131 => x"00", -- $0f2b3
          62132 => x"00", -- $0f2b4
          62133 => x"00", -- $0f2b5
          62134 => x"00", -- $0f2b6
          62135 => x"00", -- $0f2b7
          62136 => x"00", -- $0f2b8
          62137 => x"00", -- $0f2b9
          62138 => x"00", -- $0f2ba
          62139 => x"00", -- $0f2bb
          62140 => x"00", -- $0f2bc
          62141 => x"00", -- $0f2bd
          62142 => x"00", -- $0f2be
          62143 => x"00", -- $0f2bf
          62144 => x"00", -- $0f2c0
          62145 => x"00", -- $0f2c1
          62146 => x"00", -- $0f2c2
          62147 => x"00", -- $0f2c3
          62148 => x"00", -- $0f2c4
          62149 => x"00", -- $0f2c5
          62150 => x"00", -- $0f2c6
          62151 => x"00", -- $0f2c7
          62152 => x"00", -- $0f2c8
          62153 => x"00", -- $0f2c9
          62154 => x"00", -- $0f2ca
          62155 => x"00", -- $0f2cb
          62156 => x"00", -- $0f2cc
          62157 => x"00", -- $0f2cd
          62158 => x"00", -- $0f2ce
          62159 => x"00", -- $0f2cf
          62160 => x"00", -- $0f2d0
          62161 => x"00", -- $0f2d1
          62162 => x"00", -- $0f2d2
          62163 => x"00", -- $0f2d3
          62164 => x"00", -- $0f2d4
          62165 => x"00", -- $0f2d5
          62166 => x"00", -- $0f2d6
          62167 => x"00", -- $0f2d7
          62168 => x"00", -- $0f2d8
          62169 => x"00", -- $0f2d9
          62170 => x"00", -- $0f2da
          62171 => x"00", -- $0f2db
          62172 => x"00", -- $0f2dc
          62173 => x"00", -- $0f2dd
          62174 => x"00", -- $0f2de
          62175 => x"00", -- $0f2df
          62176 => x"00", -- $0f2e0
          62177 => x"00", -- $0f2e1
          62178 => x"00", -- $0f2e2
          62179 => x"00", -- $0f2e3
          62180 => x"00", -- $0f2e4
          62181 => x"00", -- $0f2e5
          62182 => x"00", -- $0f2e6
          62183 => x"00", -- $0f2e7
          62184 => x"00", -- $0f2e8
          62185 => x"00", -- $0f2e9
          62186 => x"00", -- $0f2ea
          62187 => x"00", -- $0f2eb
          62188 => x"00", -- $0f2ec
          62189 => x"00", -- $0f2ed
          62190 => x"00", -- $0f2ee
          62191 => x"00", -- $0f2ef
          62192 => x"00", -- $0f2f0
          62193 => x"00", -- $0f2f1
          62194 => x"00", -- $0f2f2
          62195 => x"00", -- $0f2f3
          62196 => x"00", -- $0f2f4
          62197 => x"00", -- $0f2f5
          62198 => x"00", -- $0f2f6
          62199 => x"00", -- $0f2f7
          62200 => x"00", -- $0f2f8
          62201 => x"00", -- $0f2f9
          62202 => x"00", -- $0f2fa
          62203 => x"00", -- $0f2fb
          62204 => x"00", -- $0f2fc
          62205 => x"00", -- $0f2fd
          62206 => x"00", -- $0f2fe
          62207 => x"00", -- $0f2ff
          62208 => x"00", -- $0f300
          62209 => x"00", -- $0f301
          62210 => x"00", -- $0f302
          62211 => x"00", -- $0f303
          62212 => x"00", -- $0f304
          62213 => x"00", -- $0f305
          62214 => x"00", -- $0f306
          62215 => x"00", -- $0f307
          62216 => x"00", -- $0f308
          62217 => x"00", -- $0f309
          62218 => x"00", -- $0f30a
          62219 => x"00", -- $0f30b
          62220 => x"00", -- $0f30c
          62221 => x"00", -- $0f30d
          62222 => x"00", -- $0f30e
          62223 => x"00", -- $0f30f
          62224 => x"00", -- $0f310
          62225 => x"00", -- $0f311
          62226 => x"00", -- $0f312
          62227 => x"00", -- $0f313
          62228 => x"00", -- $0f314
          62229 => x"00", -- $0f315
          62230 => x"00", -- $0f316
          62231 => x"00", -- $0f317
          62232 => x"00", -- $0f318
          62233 => x"00", -- $0f319
          62234 => x"00", -- $0f31a
          62235 => x"00", -- $0f31b
          62236 => x"00", -- $0f31c
          62237 => x"00", -- $0f31d
          62238 => x"00", -- $0f31e
          62239 => x"00", -- $0f31f
          62240 => x"00", -- $0f320
          62241 => x"00", -- $0f321
          62242 => x"00", -- $0f322
          62243 => x"00", -- $0f323
          62244 => x"00", -- $0f324
          62245 => x"00", -- $0f325
          62246 => x"00", -- $0f326
          62247 => x"00", -- $0f327
          62248 => x"00", -- $0f328
          62249 => x"00", -- $0f329
          62250 => x"00", -- $0f32a
          62251 => x"00", -- $0f32b
          62252 => x"00", -- $0f32c
          62253 => x"00", -- $0f32d
          62254 => x"00", -- $0f32e
          62255 => x"00", -- $0f32f
          62256 => x"00", -- $0f330
          62257 => x"00", -- $0f331
          62258 => x"00", -- $0f332
          62259 => x"00", -- $0f333
          62260 => x"00", -- $0f334
          62261 => x"00", -- $0f335
          62262 => x"00", -- $0f336
          62263 => x"00", -- $0f337
          62264 => x"00", -- $0f338
          62265 => x"00", -- $0f339
          62266 => x"00", -- $0f33a
          62267 => x"00", -- $0f33b
          62268 => x"00", -- $0f33c
          62269 => x"00", -- $0f33d
          62270 => x"00", -- $0f33e
          62271 => x"00", -- $0f33f
          62272 => x"00", -- $0f340
          62273 => x"00", -- $0f341
          62274 => x"00", -- $0f342
          62275 => x"00", -- $0f343
          62276 => x"00", -- $0f344
          62277 => x"00", -- $0f345
          62278 => x"00", -- $0f346
          62279 => x"00", -- $0f347
          62280 => x"00", -- $0f348
          62281 => x"00", -- $0f349
          62282 => x"00", -- $0f34a
          62283 => x"00", -- $0f34b
          62284 => x"00", -- $0f34c
          62285 => x"00", -- $0f34d
          62286 => x"00", -- $0f34e
          62287 => x"00", -- $0f34f
          62288 => x"00", -- $0f350
          62289 => x"00", -- $0f351
          62290 => x"00", -- $0f352
          62291 => x"00", -- $0f353
          62292 => x"00", -- $0f354
          62293 => x"00", -- $0f355
          62294 => x"00", -- $0f356
          62295 => x"00", -- $0f357
          62296 => x"00", -- $0f358
          62297 => x"00", -- $0f359
          62298 => x"00", -- $0f35a
          62299 => x"00", -- $0f35b
          62300 => x"00", -- $0f35c
          62301 => x"00", -- $0f35d
          62302 => x"00", -- $0f35e
          62303 => x"00", -- $0f35f
          62304 => x"00", -- $0f360
          62305 => x"00", -- $0f361
          62306 => x"00", -- $0f362
          62307 => x"00", -- $0f363
          62308 => x"00", -- $0f364
          62309 => x"00", -- $0f365
          62310 => x"00", -- $0f366
          62311 => x"00", -- $0f367
          62312 => x"00", -- $0f368
          62313 => x"00", -- $0f369
          62314 => x"00", -- $0f36a
          62315 => x"00", -- $0f36b
          62316 => x"00", -- $0f36c
          62317 => x"00", -- $0f36d
          62318 => x"00", -- $0f36e
          62319 => x"00", -- $0f36f
          62320 => x"00", -- $0f370
          62321 => x"00", -- $0f371
          62322 => x"00", -- $0f372
          62323 => x"00", -- $0f373
          62324 => x"00", -- $0f374
          62325 => x"00", -- $0f375
          62326 => x"00", -- $0f376
          62327 => x"00", -- $0f377
          62328 => x"00", -- $0f378
          62329 => x"00", -- $0f379
          62330 => x"00", -- $0f37a
          62331 => x"00", -- $0f37b
          62332 => x"00", -- $0f37c
          62333 => x"00", -- $0f37d
          62334 => x"00", -- $0f37e
          62335 => x"00", -- $0f37f
          62336 => x"00", -- $0f380
          62337 => x"00", -- $0f381
          62338 => x"00", -- $0f382
          62339 => x"00", -- $0f383
          62340 => x"00", -- $0f384
          62341 => x"00", -- $0f385
          62342 => x"00", -- $0f386
          62343 => x"00", -- $0f387
          62344 => x"00", -- $0f388
          62345 => x"00", -- $0f389
          62346 => x"00", -- $0f38a
          62347 => x"00", -- $0f38b
          62348 => x"00", -- $0f38c
          62349 => x"00", -- $0f38d
          62350 => x"00", -- $0f38e
          62351 => x"00", -- $0f38f
          62352 => x"00", -- $0f390
          62353 => x"00", -- $0f391
          62354 => x"00", -- $0f392
          62355 => x"00", -- $0f393
          62356 => x"00", -- $0f394
          62357 => x"00", -- $0f395
          62358 => x"00", -- $0f396
          62359 => x"00", -- $0f397
          62360 => x"00", -- $0f398
          62361 => x"00", -- $0f399
          62362 => x"00", -- $0f39a
          62363 => x"00", -- $0f39b
          62364 => x"00", -- $0f39c
          62365 => x"00", -- $0f39d
          62366 => x"00", -- $0f39e
          62367 => x"00", -- $0f39f
          62368 => x"00", -- $0f3a0
          62369 => x"00", -- $0f3a1
          62370 => x"00", -- $0f3a2
          62371 => x"00", -- $0f3a3
          62372 => x"00", -- $0f3a4
          62373 => x"00", -- $0f3a5
          62374 => x"00", -- $0f3a6
          62375 => x"00", -- $0f3a7
          62376 => x"00", -- $0f3a8
          62377 => x"00", -- $0f3a9
          62378 => x"00", -- $0f3aa
          62379 => x"00", -- $0f3ab
          62380 => x"00", -- $0f3ac
          62381 => x"00", -- $0f3ad
          62382 => x"00", -- $0f3ae
          62383 => x"00", -- $0f3af
          62384 => x"00", -- $0f3b0
          62385 => x"00", -- $0f3b1
          62386 => x"00", -- $0f3b2
          62387 => x"00", -- $0f3b3
          62388 => x"00", -- $0f3b4
          62389 => x"00", -- $0f3b5
          62390 => x"00", -- $0f3b6
          62391 => x"00", -- $0f3b7
          62392 => x"00", -- $0f3b8
          62393 => x"00", -- $0f3b9
          62394 => x"00", -- $0f3ba
          62395 => x"00", -- $0f3bb
          62396 => x"00", -- $0f3bc
          62397 => x"00", -- $0f3bd
          62398 => x"00", -- $0f3be
          62399 => x"00", -- $0f3bf
          62400 => x"00", -- $0f3c0
          62401 => x"00", -- $0f3c1
          62402 => x"00", -- $0f3c2
          62403 => x"00", -- $0f3c3
          62404 => x"00", -- $0f3c4
          62405 => x"00", -- $0f3c5
          62406 => x"00", -- $0f3c6
          62407 => x"00", -- $0f3c7
          62408 => x"00", -- $0f3c8
          62409 => x"00", -- $0f3c9
          62410 => x"00", -- $0f3ca
          62411 => x"00", -- $0f3cb
          62412 => x"00", -- $0f3cc
          62413 => x"00", -- $0f3cd
          62414 => x"00", -- $0f3ce
          62415 => x"00", -- $0f3cf
          62416 => x"00", -- $0f3d0
          62417 => x"00", -- $0f3d1
          62418 => x"00", -- $0f3d2
          62419 => x"00", -- $0f3d3
          62420 => x"00", -- $0f3d4
          62421 => x"00", -- $0f3d5
          62422 => x"00", -- $0f3d6
          62423 => x"00", -- $0f3d7
          62424 => x"00", -- $0f3d8
          62425 => x"00", -- $0f3d9
          62426 => x"00", -- $0f3da
          62427 => x"00", -- $0f3db
          62428 => x"00", -- $0f3dc
          62429 => x"00", -- $0f3dd
          62430 => x"00", -- $0f3de
          62431 => x"00", -- $0f3df
          62432 => x"00", -- $0f3e0
          62433 => x"00", -- $0f3e1
          62434 => x"00", -- $0f3e2
          62435 => x"00", -- $0f3e3
          62436 => x"00", -- $0f3e4
          62437 => x"00", -- $0f3e5
          62438 => x"00", -- $0f3e6
          62439 => x"00", -- $0f3e7
          62440 => x"00", -- $0f3e8
          62441 => x"00", -- $0f3e9
          62442 => x"00", -- $0f3ea
          62443 => x"00", -- $0f3eb
          62444 => x"00", -- $0f3ec
          62445 => x"00", -- $0f3ed
          62446 => x"00", -- $0f3ee
          62447 => x"00", -- $0f3ef
          62448 => x"00", -- $0f3f0
          62449 => x"00", -- $0f3f1
          62450 => x"00", -- $0f3f2
          62451 => x"00", -- $0f3f3
          62452 => x"00", -- $0f3f4
          62453 => x"00", -- $0f3f5
          62454 => x"00", -- $0f3f6
          62455 => x"00", -- $0f3f7
          62456 => x"00", -- $0f3f8
          62457 => x"00", -- $0f3f9
          62458 => x"00", -- $0f3fa
          62459 => x"00", -- $0f3fb
          62460 => x"00", -- $0f3fc
          62461 => x"00", -- $0f3fd
          62462 => x"00", -- $0f3fe
          62463 => x"00", -- $0f3ff
          62464 => x"00", -- $0f400
          62465 => x"00", -- $0f401
          62466 => x"00", -- $0f402
          62467 => x"00", -- $0f403
          62468 => x"00", -- $0f404
          62469 => x"00", -- $0f405
          62470 => x"00", -- $0f406
          62471 => x"00", -- $0f407
          62472 => x"00", -- $0f408
          62473 => x"00", -- $0f409
          62474 => x"00", -- $0f40a
          62475 => x"00", -- $0f40b
          62476 => x"00", -- $0f40c
          62477 => x"00", -- $0f40d
          62478 => x"00", -- $0f40e
          62479 => x"00", -- $0f40f
          62480 => x"00", -- $0f410
          62481 => x"00", -- $0f411
          62482 => x"00", -- $0f412
          62483 => x"00", -- $0f413
          62484 => x"00", -- $0f414
          62485 => x"00", -- $0f415
          62486 => x"00", -- $0f416
          62487 => x"00", -- $0f417
          62488 => x"00", -- $0f418
          62489 => x"00", -- $0f419
          62490 => x"00", -- $0f41a
          62491 => x"00", -- $0f41b
          62492 => x"00", -- $0f41c
          62493 => x"00", -- $0f41d
          62494 => x"00", -- $0f41e
          62495 => x"00", -- $0f41f
          62496 => x"00", -- $0f420
          62497 => x"00", -- $0f421
          62498 => x"00", -- $0f422
          62499 => x"00", -- $0f423
          62500 => x"00", -- $0f424
          62501 => x"00", -- $0f425
          62502 => x"00", -- $0f426
          62503 => x"00", -- $0f427
          62504 => x"00", -- $0f428
          62505 => x"00", -- $0f429
          62506 => x"00", -- $0f42a
          62507 => x"00", -- $0f42b
          62508 => x"00", -- $0f42c
          62509 => x"00", -- $0f42d
          62510 => x"00", -- $0f42e
          62511 => x"00", -- $0f42f
          62512 => x"00", -- $0f430
          62513 => x"00", -- $0f431
          62514 => x"00", -- $0f432
          62515 => x"00", -- $0f433
          62516 => x"00", -- $0f434
          62517 => x"00", -- $0f435
          62518 => x"00", -- $0f436
          62519 => x"00", -- $0f437
          62520 => x"00", -- $0f438
          62521 => x"00", -- $0f439
          62522 => x"00", -- $0f43a
          62523 => x"00", -- $0f43b
          62524 => x"00", -- $0f43c
          62525 => x"00", -- $0f43d
          62526 => x"00", -- $0f43e
          62527 => x"00", -- $0f43f
          62528 => x"00", -- $0f440
          62529 => x"00", -- $0f441
          62530 => x"00", -- $0f442
          62531 => x"00", -- $0f443
          62532 => x"00", -- $0f444
          62533 => x"00", -- $0f445
          62534 => x"00", -- $0f446
          62535 => x"00", -- $0f447
          62536 => x"00", -- $0f448
          62537 => x"00", -- $0f449
          62538 => x"00", -- $0f44a
          62539 => x"00", -- $0f44b
          62540 => x"00", -- $0f44c
          62541 => x"00", -- $0f44d
          62542 => x"00", -- $0f44e
          62543 => x"00", -- $0f44f
          62544 => x"00", -- $0f450
          62545 => x"00", -- $0f451
          62546 => x"00", -- $0f452
          62547 => x"00", -- $0f453
          62548 => x"00", -- $0f454
          62549 => x"00", -- $0f455
          62550 => x"00", -- $0f456
          62551 => x"00", -- $0f457
          62552 => x"00", -- $0f458
          62553 => x"00", -- $0f459
          62554 => x"00", -- $0f45a
          62555 => x"00", -- $0f45b
          62556 => x"00", -- $0f45c
          62557 => x"00", -- $0f45d
          62558 => x"00", -- $0f45e
          62559 => x"00", -- $0f45f
          62560 => x"00", -- $0f460
          62561 => x"00", -- $0f461
          62562 => x"00", -- $0f462
          62563 => x"00", -- $0f463
          62564 => x"00", -- $0f464
          62565 => x"00", -- $0f465
          62566 => x"00", -- $0f466
          62567 => x"00", -- $0f467
          62568 => x"00", -- $0f468
          62569 => x"00", -- $0f469
          62570 => x"00", -- $0f46a
          62571 => x"00", -- $0f46b
          62572 => x"00", -- $0f46c
          62573 => x"00", -- $0f46d
          62574 => x"00", -- $0f46e
          62575 => x"00", -- $0f46f
          62576 => x"00", -- $0f470
          62577 => x"00", -- $0f471
          62578 => x"00", -- $0f472
          62579 => x"00", -- $0f473
          62580 => x"00", -- $0f474
          62581 => x"00", -- $0f475
          62582 => x"00", -- $0f476
          62583 => x"00", -- $0f477
          62584 => x"00", -- $0f478
          62585 => x"00", -- $0f479
          62586 => x"00", -- $0f47a
          62587 => x"00", -- $0f47b
          62588 => x"00", -- $0f47c
          62589 => x"00", -- $0f47d
          62590 => x"00", -- $0f47e
          62591 => x"00", -- $0f47f
          62592 => x"00", -- $0f480
          62593 => x"00", -- $0f481
          62594 => x"00", -- $0f482
          62595 => x"00", -- $0f483
          62596 => x"00", -- $0f484
          62597 => x"00", -- $0f485
          62598 => x"00", -- $0f486
          62599 => x"00", -- $0f487
          62600 => x"00", -- $0f488
          62601 => x"00", -- $0f489
          62602 => x"00", -- $0f48a
          62603 => x"00", -- $0f48b
          62604 => x"00", -- $0f48c
          62605 => x"00", -- $0f48d
          62606 => x"00", -- $0f48e
          62607 => x"00", -- $0f48f
          62608 => x"00", -- $0f490
          62609 => x"00", -- $0f491
          62610 => x"00", -- $0f492
          62611 => x"00", -- $0f493
          62612 => x"00", -- $0f494
          62613 => x"00", -- $0f495
          62614 => x"00", -- $0f496
          62615 => x"00", -- $0f497
          62616 => x"00", -- $0f498
          62617 => x"00", -- $0f499
          62618 => x"00", -- $0f49a
          62619 => x"00", -- $0f49b
          62620 => x"00", -- $0f49c
          62621 => x"00", -- $0f49d
          62622 => x"00", -- $0f49e
          62623 => x"00", -- $0f49f
          62624 => x"00", -- $0f4a0
          62625 => x"00", -- $0f4a1
          62626 => x"00", -- $0f4a2
          62627 => x"00", -- $0f4a3
          62628 => x"00", -- $0f4a4
          62629 => x"00", -- $0f4a5
          62630 => x"00", -- $0f4a6
          62631 => x"00", -- $0f4a7
          62632 => x"00", -- $0f4a8
          62633 => x"00", -- $0f4a9
          62634 => x"00", -- $0f4aa
          62635 => x"00", -- $0f4ab
          62636 => x"00", -- $0f4ac
          62637 => x"00", -- $0f4ad
          62638 => x"00", -- $0f4ae
          62639 => x"00", -- $0f4af
          62640 => x"00", -- $0f4b0
          62641 => x"00", -- $0f4b1
          62642 => x"00", -- $0f4b2
          62643 => x"00", -- $0f4b3
          62644 => x"00", -- $0f4b4
          62645 => x"00", -- $0f4b5
          62646 => x"00", -- $0f4b6
          62647 => x"00", -- $0f4b7
          62648 => x"00", -- $0f4b8
          62649 => x"00", -- $0f4b9
          62650 => x"00", -- $0f4ba
          62651 => x"00", -- $0f4bb
          62652 => x"00", -- $0f4bc
          62653 => x"00", -- $0f4bd
          62654 => x"00", -- $0f4be
          62655 => x"00", -- $0f4bf
          62656 => x"00", -- $0f4c0
          62657 => x"00", -- $0f4c1
          62658 => x"00", -- $0f4c2
          62659 => x"00", -- $0f4c3
          62660 => x"00", -- $0f4c4
          62661 => x"00", -- $0f4c5
          62662 => x"00", -- $0f4c6
          62663 => x"00", -- $0f4c7
          62664 => x"00", -- $0f4c8
          62665 => x"00", -- $0f4c9
          62666 => x"00", -- $0f4ca
          62667 => x"00", -- $0f4cb
          62668 => x"00", -- $0f4cc
          62669 => x"00", -- $0f4cd
          62670 => x"00", -- $0f4ce
          62671 => x"00", -- $0f4cf
          62672 => x"00", -- $0f4d0
          62673 => x"00", -- $0f4d1
          62674 => x"00", -- $0f4d2
          62675 => x"00", -- $0f4d3
          62676 => x"00", -- $0f4d4
          62677 => x"00", -- $0f4d5
          62678 => x"00", -- $0f4d6
          62679 => x"00", -- $0f4d7
          62680 => x"00", -- $0f4d8
          62681 => x"00", -- $0f4d9
          62682 => x"00", -- $0f4da
          62683 => x"00", -- $0f4db
          62684 => x"00", -- $0f4dc
          62685 => x"00", -- $0f4dd
          62686 => x"00", -- $0f4de
          62687 => x"00", -- $0f4df
          62688 => x"00", -- $0f4e0
          62689 => x"00", -- $0f4e1
          62690 => x"00", -- $0f4e2
          62691 => x"00", -- $0f4e3
          62692 => x"00", -- $0f4e4
          62693 => x"00", -- $0f4e5
          62694 => x"00", -- $0f4e6
          62695 => x"00", -- $0f4e7
          62696 => x"00", -- $0f4e8
          62697 => x"00", -- $0f4e9
          62698 => x"00", -- $0f4ea
          62699 => x"00", -- $0f4eb
          62700 => x"00", -- $0f4ec
          62701 => x"00", -- $0f4ed
          62702 => x"00", -- $0f4ee
          62703 => x"00", -- $0f4ef
          62704 => x"00", -- $0f4f0
          62705 => x"00", -- $0f4f1
          62706 => x"00", -- $0f4f2
          62707 => x"00", -- $0f4f3
          62708 => x"00", -- $0f4f4
          62709 => x"00", -- $0f4f5
          62710 => x"00", -- $0f4f6
          62711 => x"00", -- $0f4f7
          62712 => x"00", -- $0f4f8
          62713 => x"00", -- $0f4f9
          62714 => x"00", -- $0f4fa
          62715 => x"00", -- $0f4fb
          62716 => x"00", -- $0f4fc
          62717 => x"00", -- $0f4fd
          62718 => x"00", -- $0f4fe
          62719 => x"00", -- $0f4ff
          62720 => x"00", -- $0f500
          62721 => x"00", -- $0f501
          62722 => x"00", -- $0f502
          62723 => x"00", -- $0f503
          62724 => x"00", -- $0f504
          62725 => x"00", -- $0f505
          62726 => x"00", -- $0f506
          62727 => x"00", -- $0f507
          62728 => x"00", -- $0f508
          62729 => x"00", -- $0f509
          62730 => x"00", -- $0f50a
          62731 => x"00", -- $0f50b
          62732 => x"00", -- $0f50c
          62733 => x"00", -- $0f50d
          62734 => x"00", -- $0f50e
          62735 => x"00", -- $0f50f
          62736 => x"00", -- $0f510
          62737 => x"00", -- $0f511
          62738 => x"00", -- $0f512
          62739 => x"00", -- $0f513
          62740 => x"00", -- $0f514
          62741 => x"00", -- $0f515
          62742 => x"00", -- $0f516
          62743 => x"00", -- $0f517
          62744 => x"00", -- $0f518
          62745 => x"00", -- $0f519
          62746 => x"00", -- $0f51a
          62747 => x"00", -- $0f51b
          62748 => x"00", -- $0f51c
          62749 => x"00", -- $0f51d
          62750 => x"00", -- $0f51e
          62751 => x"00", -- $0f51f
          62752 => x"00", -- $0f520
          62753 => x"00", -- $0f521
          62754 => x"00", -- $0f522
          62755 => x"00", -- $0f523
          62756 => x"00", -- $0f524
          62757 => x"00", -- $0f525
          62758 => x"00", -- $0f526
          62759 => x"00", -- $0f527
          62760 => x"00", -- $0f528
          62761 => x"00", -- $0f529
          62762 => x"00", -- $0f52a
          62763 => x"00", -- $0f52b
          62764 => x"00", -- $0f52c
          62765 => x"00", -- $0f52d
          62766 => x"00", -- $0f52e
          62767 => x"00", -- $0f52f
          62768 => x"00", -- $0f530
          62769 => x"00", -- $0f531
          62770 => x"00", -- $0f532
          62771 => x"00", -- $0f533
          62772 => x"00", -- $0f534
          62773 => x"00", -- $0f535
          62774 => x"00", -- $0f536
          62775 => x"00", -- $0f537
          62776 => x"00", -- $0f538
          62777 => x"00", -- $0f539
          62778 => x"00", -- $0f53a
          62779 => x"00", -- $0f53b
          62780 => x"00", -- $0f53c
          62781 => x"00", -- $0f53d
          62782 => x"00", -- $0f53e
          62783 => x"00", -- $0f53f
          62784 => x"00", -- $0f540
          62785 => x"00", -- $0f541
          62786 => x"00", -- $0f542
          62787 => x"00", -- $0f543
          62788 => x"00", -- $0f544
          62789 => x"00", -- $0f545
          62790 => x"00", -- $0f546
          62791 => x"00", -- $0f547
          62792 => x"00", -- $0f548
          62793 => x"00", -- $0f549
          62794 => x"00", -- $0f54a
          62795 => x"00", -- $0f54b
          62796 => x"00", -- $0f54c
          62797 => x"00", -- $0f54d
          62798 => x"00", -- $0f54e
          62799 => x"00", -- $0f54f
          62800 => x"00", -- $0f550
          62801 => x"00", -- $0f551
          62802 => x"00", -- $0f552
          62803 => x"00", -- $0f553
          62804 => x"00", -- $0f554
          62805 => x"00", -- $0f555
          62806 => x"00", -- $0f556
          62807 => x"00", -- $0f557
          62808 => x"00", -- $0f558
          62809 => x"00", -- $0f559
          62810 => x"00", -- $0f55a
          62811 => x"00", -- $0f55b
          62812 => x"00", -- $0f55c
          62813 => x"00", -- $0f55d
          62814 => x"00", -- $0f55e
          62815 => x"00", -- $0f55f
          62816 => x"00", -- $0f560
          62817 => x"00", -- $0f561
          62818 => x"00", -- $0f562
          62819 => x"00", -- $0f563
          62820 => x"00", -- $0f564
          62821 => x"00", -- $0f565
          62822 => x"00", -- $0f566
          62823 => x"00", -- $0f567
          62824 => x"00", -- $0f568
          62825 => x"00", -- $0f569
          62826 => x"00", -- $0f56a
          62827 => x"00", -- $0f56b
          62828 => x"00", -- $0f56c
          62829 => x"00", -- $0f56d
          62830 => x"00", -- $0f56e
          62831 => x"00", -- $0f56f
          62832 => x"00", -- $0f570
          62833 => x"00", -- $0f571
          62834 => x"00", -- $0f572
          62835 => x"00", -- $0f573
          62836 => x"00", -- $0f574
          62837 => x"00", -- $0f575
          62838 => x"00", -- $0f576
          62839 => x"00", -- $0f577
          62840 => x"00", -- $0f578
          62841 => x"00", -- $0f579
          62842 => x"00", -- $0f57a
          62843 => x"00", -- $0f57b
          62844 => x"00", -- $0f57c
          62845 => x"00", -- $0f57d
          62846 => x"00", -- $0f57e
          62847 => x"00", -- $0f57f
          62848 => x"00", -- $0f580
          62849 => x"00", -- $0f581
          62850 => x"00", -- $0f582
          62851 => x"00", -- $0f583
          62852 => x"00", -- $0f584
          62853 => x"00", -- $0f585
          62854 => x"00", -- $0f586
          62855 => x"00", -- $0f587
          62856 => x"00", -- $0f588
          62857 => x"00", -- $0f589
          62858 => x"00", -- $0f58a
          62859 => x"00", -- $0f58b
          62860 => x"00", -- $0f58c
          62861 => x"00", -- $0f58d
          62862 => x"00", -- $0f58e
          62863 => x"00", -- $0f58f
          62864 => x"00", -- $0f590
          62865 => x"00", -- $0f591
          62866 => x"00", -- $0f592
          62867 => x"00", -- $0f593
          62868 => x"00", -- $0f594
          62869 => x"00", -- $0f595
          62870 => x"00", -- $0f596
          62871 => x"00", -- $0f597
          62872 => x"00", -- $0f598
          62873 => x"00", -- $0f599
          62874 => x"00", -- $0f59a
          62875 => x"00", -- $0f59b
          62876 => x"00", -- $0f59c
          62877 => x"00", -- $0f59d
          62878 => x"00", -- $0f59e
          62879 => x"00", -- $0f59f
          62880 => x"00", -- $0f5a0
          62881 => x"00", -- $0f5a1
          62882 => x"00", -- $0f5a2
          62883 => x"00", -- $0f5a3
          62884 => x"00", -- $0f5a4
          62885 => x"00", -- $0f5a5
          62886 => x"00", -- $0f5a6
          62887 => x"00", -- $0f5a7
          62888 => x"00", -- $0f5a8
          62889 => x"00", -- $0f5a9
          62890 => x"00", -- $0f5aa
          62891 => x"00", -- $0f5ab
          62892 => x"00", -- $0f5ac
          62893 => x"00", -- $0f5ad
          62894 => x"00", -- $0f5ae
          62895 => x"00", -- $0f5af
          62896 => x"00", -- $0f5b0
          62897 => x"00", -- $0f5b1
          62898 => x"00", -- $0f5b2
          62899 => x"00", -- $0f5b3
          62900 => x"00", -- $0f5b4
          62901 => x"00", -- $0f5b5
          62902 => x"00", -- $0f5b6
          62903 => x"00", -- $0f5b7
          62904 => x"00", -- $0f5b8
          62905 => x"00", -- $0f5b9
          62906 => x"00", -- $0f5ba
          62907 => x"00", -- $0f5bb
          62908 => x"00", -- $0f5bc
          62909 => x"00", -- $0f5bd
          62910 => x"00", -- $0f5be
          62911 => x"00", -- $0f5bf
          62912 => x"00", -- $0f5c0
          62913 => x"00", -- $0f5c1
          62914 => x"00", -- $0f5c2
          62915 => x"00", -- $0f5c3
          62916 => x"00", -- $0f5c4
          62917 => x"00", -- $0f5c5
          62918 => x"00", -- $0f5c6
          62919 => x"00", -- $0f5c7
          62920 => x"00", -- $0f5c8
          62921 => x"00", -- $0f5c9
          62922 => x"00", -- $0f5ca
          62923 => x"00", -- $0f5cb
          62924 => x"00", -- $0f5cc
          62925 => x"00", -- $0f5cd
          62926 => x"00", -- $0f5ce
          62927 => x"00", -- $0f5cf
          62928 => x"00", -- $0f5d0
          62929 => x"00", -- $0f5d1
          62930 => x"00", -- $0f5d2
          62931 => x"00", -- $0f5d3
          62932 => x"00", -- $0f5d4
          62933 => x"00", -- $0f5d5
          62934 => x"00", -- $0f5d6
          62935 => x"00", -- $0f5d7
          62936 => x"00", -- $0f5d8
          62937 => x"00", -- $0f5d9
          62938 => x"00", -- $0f5da
          62939 => x"00", -- $0f5db
          62940 => x"00", -- $0f5dc
          62941 => x"00", -- $0f5dd
          62942 => x"00", -- $0f5de
          62943 => x"00", -- $0f5df
          62944 => x"00", -- $0f5e0
          62945 => x"00", -- $0f5e1
          62946 => x"00", -- $0f5e2
          62947 => x"00", -- $0f5e3
          62948 => x"00", -- $0f5e4
          62949 => x"00", -- $0f5e5
          62950 => x"00", -- $0f5e6
          62951 => x"00", -- $0f5e7
          62952 => x"00", -- $0f5e8
          62953 => x"00", -- $0f5e9
          62954 => x"00", -- $0f5ea
          62955 => x"00", -- $0f5eb
          62956 => x"00", -- $0f5ec
          62957 => x"00", -- $0f5ed
          62958 => x"00", -- $0f5ee
          62959 => x"00", -- $0f5ef
          62960 => x"00", -- $0f5f0
          62961 => x"00", -- $0f5f1
          62962 => x"00", -- $0f5f2
          62963 => x"00", -- $0f5f3
          62964 => x"00", -- $0f5f4
          62965 => x"00", -- $0f5f5
          62966 => x"00", -- $0f5f6
          62967 => x"00", -- $0f5f7
          62968 => x"00", -- $0f5f8
          62969 => x"00", -- $0f5f9
          62970 => x"00", -- $0f5fa
          62971 => x"00", -- $0f5fb
          62972 => x"00", -- $0f5fc
          62973 => x"00", -- $0f5fd
          62974 => x"00", -- $0f5fe
          62975 => x"00", -- $0f5ff
          62976 => x"00", -- $0f600
          62977 => x"00", -- $0f601
          62978 => x"00", -- $0f602
          62979 => x"00", -- $0f603
          62980 => x"00", -- $0f604
          62981 => x"00", -- $0f605
          62982 => x"00", -- $0f606
          62983 => x"00", -- $0f607
          62984 => x"00", -- $0f608
          62985 => x"00", -- $0f609
          62986 => x"00", -- $0f60a
          62987 => x"00", -- $0f60b
          62988 => x"00", -- $0f60c
          62989 => x"00", -- $0f60d
          62990 => x"00", -- $0f60e
          62991 => x"00", -- $0f60f
          62992 => x"00", -- $0f610
          62993 => x"00", -- $0f611
          62994 => x"00", -- $0f612
          62995 => x"00", -- $0f613
          62996 => x"00", -- $0f614
          62997 => x"00", -- $0f615
          62998 => x"00", -- $0f616
          62999 => x"00", -- $0f617
          63000 => x"00", -- $0f618
          63001 => x"00", -- $0f619
          63002 => x"00", -- $0f61a
          63003 => x"00", -- $0f61b
          63004 => x"00", -- $0f61c
          63005 => x"00", -- $0f61d
          63006 => x"00", -- $0f61e
          63007 => x"00", -- $0f61f
          63008 => x"00", -- $0f620
          63009 => x"00", -- $0f621
          63010 => x"00", -- $0f622
          63011 => x"00", -- $0f623
          63012 => x"00", -- $0f624
          63013 => x"00", -- $0f625
          63014 => x"00", -- $0f626
          63015 => x"00", -- $0f627
          63016 => x"00", -- $0f628
          63017 => x"00", -- $0f629
          63018 => x"00", -- $0f62a
          63019 => x"00", -- $0f62b
          63020 => x"00", -- $0f62c
          63021 => x"00", -- $0f62d
          63022 => x"00", -- $0f62e
          63023 => x"00", -- $0f62f
          63024 => x"00", -- $0f630
          63025 => x"00", -- $0f631
          63026 => x"00", -- $0f632
          63027 => x"00", -- $0f633
          63028 => x"00", -- $0f634
          63029 => x"00", -- $0f635
          63030 => x"00", -- $0f636
          63031 => x"00", -- $0f637
          63032 => x"00", -- $0f638
          63033 => x"00", -- $0f639
          63034 => x"00", -- $0f63a
          63035 => x"00", -- $0f63b
          63036 => x"00", -- $0f63c
          63037 => x"00", -- $0f63d
          63038 => x"00", -- $0f63e
          63039 => x"00", -- $0f63f
          63040 => x"00", -- $0f640
          63041 => x"00", -- $0f641
          63042 => x"00", -- $0f642
          63043 => x"00", -- $0f643
          63044 => x"00", -- $0f644
          63045 => x"00", -- $0f645
          63046 => x"00", -- $0f646
          63047 => x"00", -- $0f647
          63048 => x"00", -- $0f648
          63049 => x"00", -- $0f649
          63050 => x"00", -- $0f64a
          63051 => x"00", -- $0f64b
          63052 => x"00", -- $0f64c
          63053 => x"00", -- $0f64d
          63054 => x"00", -- $0f64e
          63055 => x"00", -- $0f64f
          63056 => x"00", -- $0f650
          63057 => x"00", -- $0f651
          63058 => x"00", -- $0f652
          63059 => x"00", -- $0f653
          63060 => x"00", -- $0f654
          63061 => x"00", -- $0f655
          63062 => x"00", -- $0f656
          63063 => x"00", -- $0f657
          63064 => x"00", -- $0f658
          63065 => x"00", -- $0f659
          63066 => x"00", -- $0f65a
          63067 => x"00", -- $0f65b
          63068 => x"00", -- $0f65c
          63069 => x"00", -- $0f65d
          63070 => x"00", -- $0f65e
          63071 => x"00", -- $0f65f
          63072 => x"00", -- $0f660
          63073 => x"00", -- $0f661
          63074 => x"00", -- $0f662
          63075 => x"00", -- $0f663
          63076 => x"00", -- $0f664
          63077 => x"00", -- $0f665
          63078 => x"00", -- $0f666
          63079 => x"00", -- $0f667
          63080 => x"00", -- $0f668
          63081 => x"00", -- $0f669
          63082 => x"00", -- $0f66a
          63083 => x"00", -- $0f66b
          63084 => x"00", -- $0f66c
          63085 => x"00", -- $0f66d
          63086 => x"00", -- $0f66e
          63087 => x"00", -- $0f66f
          63088 => x"00", -- $0f670
          63089 => x"00", -- $0f671
          63090 => x"00", -- $0f672
          63091 => x"00", -- $0f673
          63092 => x"00", -- $0f674
          63093 => x"00", -- $0f675
          63094 => x"00", -- $0f676
          63095 => x"00", -- $0f677
          63096 => x"00", -- $0f678
          63097 => x"00", -- $0f679
          63098 => x"00", -- $0f67a
          63099 => x"00", -- $0f67b
          63100 => x"00", -- $0f67c
          63101 => x"00", -- $0f67d
          63102 => x"00", -- $0f67e
          63103 => x"00", -- $0f67f
          63104 => x"00", -- $0f680
          63105 => x"00", -- $0f681
          63106 => x"00", -- $0f682
          63107 => x"00", -- $0f683
          63108 => x"00", -- $0f684
          63109 => x"00", -- $0f685
          63110 => x"00", -- $0f686
          63111 => x"00", -- $0f687
          63112 => x"00", -- $0f688
          63113 => x"00", -- $0f689
          63114 => x"00", -- $0f68a
          63115 => x"00", -- $0f68b
          63116 => x"00", -- $0f68c
          63117 => x"00", -- $0f68d
          63118 => x"00", -- $0f68e
          63119 => x"00", -- $0f68f
          63120 => x"00", -- $0f690
          63121 => x"00", -- $0f691
          63122 => x"00", -- $0f692
          63123 => x"00", -- $0f693
          63124 => x"00", -- $0f694
          63125 => x"00", -- $0f695
          63126 => x"00", -- $0f696
          63127 => x"00", -- $0f697
          63128 => x"00", -- $0f698
          63129 => x"00", -- $0f699
          63130 => x"00", -- $0f69a
          63131 => x"00", -- $0f69b
          63132 => x"00", -- $0f69c
          63133 => x"00", -- $0f69d
          63134 => x"00", -- $0f69e
          63135 => x"00", -- $0f69f
          63136 => x"00", -- $0f6a0
          63137 => x"00", -- $0f6a1
          63138 => x"00", -- $0f6a2
          63139 => x"00", -- $0f6a3
          63140 => x"00", -- $0f6a4
          63141 => x"00", -- $0f6a5
          63142 => x"00", -- $0f6a6
          63143 => x"00", -- $0f6a7
          63144 => x"00", -- $0f6a8
          63145 => x"00", -- $0f6a9
          63146 => x"00", -- $0f6aa
          63147 => x"00", -- $0f6ab
          63148 => x"00", -- $0f6ac
          63149 => x"00", -- $0f6ad
          63150 => x"00", -- $0f6ae
          63151 => x"00", -- $0f6af
          63152 => x"00", -- $0f6b0
          63153 => x"00", -- $0f6b1
          63154 => x"00", -- $0f6b2
          63155 => x"00", -- $0f6b3
          63156 => x"00", -- $0f6b4
          63157 => x"00", -- $0f6b5
          63158 => x"00", -- $0f6b6
          63159 => x"00", -- $0f6b7
          63160 => x"00", -- $0f6b8
          63161 => x"00", -- $0f6b9
          63162 => x"00", -- $0f6ba
          63163 => x"00", -- $0f6bb
          63164 => x"00", -- $0f6bc
          63165 => x"00", -- $0f6bd
          63166 => x"00", -- $0f6be
          63167 => x"00", -- $0f6bf
          63168 => x"00", -- $0f6c0
          63169 => x"00", -- $0f6c1
          63170 => x"00", -- $0f6c2
          63171 => x"00", -- $0f6c3
          63172 => x"00", -- $0f6c4
          63173 => x"00", -- $0f6c5
          63174 => x"00", -- $0f6c6
          63175 => x"00", -- $0f6c7
          63176 => x"00", -- $0f6c8
          63177 => x"00", -- $0f6c9
          63178 => x"00", -- $0f6ca
          63179 => x"00", -- $0f6cb
          63180 => x"00", -- $0f6cc
          63181 => x"00", -- $0f6cd
          63182 => x"00", -- $0f6ce
          63183 => x"00", -- $0f6cf
          63184 => x"00", -- $0f6d0
          63185 => x"00", -- $0f6d1
          63186 => x"00", -- $0f6d2
          63187 => x"00", -- $0f6d3
          63188 => x"00", -- $0f6d4
          63189 => x"00", -- $0f6d5
          63190 => x"00", -- $0f6d6
          63191 => x"00", -- $0f6d7
          63192 => x"00", -- $0f6d8
          63193 => x"00", -- $0f6d9
          63194 => x"00", -- $0f6da
          63195 => x"00", -- $0f6db
          63196 => x"00", -- $0f6dc
          63197 => x"00", -- $0f6dd
          63198 => x"00", -- $0f6de
          63199 => x"00", -- $0f6df
          63200 => x"00", -- $0f6e0
          63201 => x"00", -- $0f6e1
          63202 => x"00", -- $0f6e2
          63203 => x"00", -- $0f6e3
          63204 => x"00", -- $0f6e4
          63205 => x"00", -- $0f6e5
          63206 => x"00", -- $0f6e6
          63207 => x"00", -- $0f6e7
          63208 => x"00", -- $0f6e8
          63209 => x"00", -- $0f6e9
          63210 => x"00", -- $0f6ea
          63211 => x"00", -- $0f6eb
          63212 => x"00", -- $0f6ec
          63213 => x"00", -- $0f6ed
          63214 => x"00", -- $0f6ee
          63215 => x"00", -- $0f6ef
          63216 => x"00", -- $0f6f0
          63217 => x"00", -- $0f6f1
          63218 => x"00", -- $0f6f2
          63219 => x"00", -- $0f6f3
          63220 => x"00", -- $0f6f4
          63221 => x"00", -- $0f6f5
          63222 => x"00", -- $0f6f6
          63223 => x"00", -- $0f6f7
          63224 => x"00", -- $0f6f8
          63225 => x"00", -- $0f6f9
          63226 => x"00", -- $0f6fa
          63227 => x"00", -- $0f6fb
          63228 => x"00", -- $0f6fc
          63229 => x"00", -- $0f6fd
          63230 => x"00", -- $0f6fe
          63231 => x"00", -- $0f6ff
          63232 => x"00", -- $0f700
          63233 => x"00", -- $0f701
          63234 => x"00", -- $0f702
          63235 => x"00", -- $0f703
          63236 => x"00", -- $0f704
          63237 => x"00", -- $0f705
          63238 => x"00", -- $0f706
          63239 => x"00", -- $0f707
          63240 => x"00", -- $0f708
          63241 => x"00", -- $0f709
          63242 => x"00", -- $0f70a
          63243 => x"00", -- $0f70b
          63244 => x"00", -- $0f70c
          63245 => x"00", -- $0f70d
          63246 => x"00", -- $0f70e
          63247 => x"00", -- $0f70f
          63248 => x"00", -- $0f710
          63249 => x"00", -- $0f711
          63250 => x"00", -- $0f712
          63251 => x"00", -- $0f713
          63252 => x"00", -- $0f714
          63253 => x"00", -- $0f715
          63254 => x"00", -- $0f716
          63255 => x"00", -- $0f717
          63256 => x"00", -- $0f718
          63257 => x"00", -- $0f719
          63258 => x"00", -- $0f71a
          63259 => x"00", -- $0f71b
          63260 => x"00", -- $0f71c
          63261 => x"00", -- $0f71d
          63262 => x"00", -- $0f71e
          63263 => x"00", -- $0f71f
          63264 => x"00", -- $0f720
          63265 => x"00", -- $0f721
          63266 => x"00", -- $0f722
          63267 => x"00", -- $0f723
          63268 => x"00", -- $0f724
          63269 => x"00", -- $0f725
          63270 => x"00", -- $0f726
          63271 => x"00", -- $0f727
          63272 => x"00", -- $0f728
          63273 => x"00", -- $0f729
          63274 => x"00", -- $0f72a
          63275 => x"00", -- $0f72b
          63276 => x"00", -- $0f72c
          63277 => x"00", -- $0f72d
          63278 => x"00", -- $0f72e
          63279 => x"00", -- $0f72f
          63280 => x"00", -- $0f730
          63281 => x"00", -- $0f731
          63282 => x"00", -- $0f732
          63283 => x"00", -- $0f733
          63284 => x"00", -- $0f734
          63285 => x"00", -- $0f735
          63286 => x"00", -- $0f736
          63287 => x"00", -- $0f737
          63288 => x"00", -- $0f738
          63289 => x"00", -- $0f739
          63290 => x"00", -- $0f73a
          63291 => x"00", -- $0f73b
          63292 => x"00", -- $0f73c
          63293 => x"00", -- $0f73d
          63294 => x"00", -- $0f73e
          63295 => x"00", -- $0f73f
          63296 => x"00", -- $0f740
          63297 => x"00", -- $0f741
          63298 => x"00", -- $0f742
          63299 => x"00", -- $0f743
          63300 => x"00", -- $0f744
          63301 => x"00", -- $0f745
          63302 => x"00", -- $0f746
          63303 => x"00", -- $0f747
          63304 => x"00", -- $0f748
          63305 => x"00", -- $0f749
          63306 => x"00", -- $0f74a
          63307 => x"00", -- $0f74b
          63308 => x"00", -- $0f74c
          63309 => x"00", -- $0f74d
          63310 => x"00", -- $0f74e
          63311 => x"00", -- $0f74f
          63312 => x"00", -- $0f750
          63313 => x"00", -- $0f751
          63314 => x"00", -- $0f752
          63315 => x"00", -- $0f753
          63316 => x"00", -- $0f754
          63317 => x"00", -- $0f755
          63318 => x"00", -- $0f756
          63319 => x"00", -- $0f757
          63320 => x"00", -- $0f758
          63321 => x"00", -- $0f759
          63322 => x"00", -- $0f75a
          63323 => x"00", -- $0f75b
          63324 => x"00", -- $0f75c
          63325 => x"00", -- $0f75d
          63326 => x"00", -- $0f75e
          63327 => x"00", -- $0f75f
          63328 => x"00", -- $0f760
          63329 => x"00", -- $0f761
          63330 => x"00", -- $0f762
          63331 => x"00", -- $0f763
          63332 => x"00", -- $0f764
          63333 => x"00", -- $0f765
          63334 => x"00", -- $0f766
          63335 => x"00", -- $0f767
          63336 => x"00", -- $0f768
          63337 => x"00", -- $0f769
          63338 => x"00", -- $0f76a
          63339 => x"00", -- $0f76b
          63340 => x"00", -- $0f76c
          63341 => x"00", -- $0f76d
          63342 => x"00", -- $0f76e
          63343 => x"00", -- $0f76f
          63344 => x"00", -- $0f770
          63345 => x"00", -- $0f771
          63346 => x"00", -- $0f772
          63347 => x"00", -- $0f773
          63348 => x"00", -- $0f774
          63349 => x"00", -- $0f775
          63350 => x"00", -- $0f776
          63351 => x"00", -- $0f777
          63352 => x"00", -- $0f778
          63353 => x"00", -- $0f779
          63354 => x"00", -- $0f77a
          63355 => x"00", -- $0f77b
          63356 => x"00", -- $0f77c
          63357 => x"00", -- $0f77d
          63358 => x"00", -- $0f77e
          63359 => x"00", -- $0f77f
          63360 => x"00", -- $0f780
          63361 => x"00", -- $0f781
          63362 => x"00", -- $0f782
          63363 => x"00", -- $0f783
          63364 => x"00", -- $0f784
          63365 => x"00", -- $0f785
          63366 => x"00", -- $0f786
          63367 => x"00", -- $0f787
          63368 => x"00", -- $0f788
          63369 => x"00", -- $0f789
          63370 => x"00", -- $0f78a
          63371 => x"00", -- $0f78b
          63372 => x"00", -- $0f78c
          63373 => x"00", -- $0f78d
          63374 => x"00", -- $0f78e
          63375 => x"00", -- $0f78f
          63376 => x"00", -- $0f790
          63377 => x"00", -- $0f791
          63378 => x"00", -- $0f792
          63379 => x"00", -- $0f793
          63380 => x"00", -- $0f794
          63381 => x"00", -- $0f795
          63382 => x"00", -- $0f796
          63383 => x"00", -- $0f797
          63384 => x"00", -- $0f798
          63385 => x"00", -- $0f799
          63386 => x"00", -- $0f79a
          63387 => x"00", -- $0f79b
          63388 => x"00", -- $0f79c
          63389 => x"00", -- $0f79d
          63390 => x"00", -- $0f79e
          63391 => x"00", -- $0f79f
          63392 => x"00", -- $0f7a0
          63393 => x"00", -- $0f7a1
          63394 => x"00", -- $0f7a2
          63395 => x"00", -- $0f7a3
          63396 => x"00", -- $0f7a4
          63397 => x"00", -- $0f7a5
          63398 => x"00", -- $0f7a6
          63399 => x"00", -- $0f7a7
          63400 => x"00", -- $0f7a8
          63401 => x"00", -- $0f7a9
          63402 => x"00", -- $0f7aa
          63403 => x"00", -- $0f7ab
          63404 => x"00", -- $0f7ac
          63405 => x"00", -- $0f7ad
          63406 => x"00", -- $0f7ae
          63407 => x"00", -- $0f7af
          63408 => x"00", -- $0f7b0
          63409 => x"00", -- $0f7b1
          63410 => x"00", -- $0f7b2
          63411 => x"00", -- $0f7b3
          63412 => x"00", -- $0f7b4
          63413 => x"00", -- $0f7b5
          63414 => x"00", -- $0f7b6
          63415 => x"00", -- $0f7b7
          63416 => x"00", -- $0f7b8
          63417 => x"00", -- $0f7b9
          63418 => x"00", -- $0f7ba
          63419 => x"00", -- $0f7bb
          63420 => x"00", -- $0f7bc
          63421 => x"00", -- $0f7bd
          63422 => x"00", -- $0f7be
          63423 => x"00", -- $0f7bf
          63424 => x"00", -- $0f7c0
          63425 => x"00", -- $0f7c1
          63426 => x"00", -- $0f7c2
          63427 => x"00", -- $0f7c3
          63428 => x"00", -- $0f7c4
          63429 => x"00", -- $0f7c5
          63430 => x"00", -- $0f7c6
          63431 => x"00", -- $0f7c7
          63432 => x"00", -- $0f7c8
          63433 => x"00", -- $0f7c9
          63434 => x"00", -- $0f7ca
          63435 => x"00", -- $0f7cb
          63436 => x"00", -- $0f7cc
          63437 => x"00", -- $0f7cd
          63438 => x"00", -- $0f7ce
          63439 => x"00", -- $0f7cf
          63440 => x"00", -- $0f7d0
          63441 => x"00", -- $0f7d1
          63442 => x"00", -- $0f7d2
          63443 => x"00", -- $0f7d3
          63444 => x"00", -- $0f7d4
          63445 => x"00", -- $0f7d5
          63446 => x"00", -- $0f7d6
          63447 => x"00", -- $0f7d7
          63448 => x"00", -- $0f7d8
          63449 => x"00", -- $0f7d9
          63450 => x"00", -- $0f7da
          63451 => x"00", -- $0f7db
          63452 => x"00", -- $0f7dc
          63453 => x"00", -- $0f7dd
          63454 => x"00", -- $0f7de
          63455 => x"00", -- $0f7df
          63456 => x"00", -- $0f7e0
          63457 => x"00", -- $0f7e1
          63458 => x"00", -- $0f7e2
          63459 => x"00", -- $0f7e3
          63460 => x"00", -- $0f7e4
          63461 => x"00", -- $0f7e5
          63462 => x"00", -- $0f7e6
          63463 => x"00", -- $0f7e7
          63464 => x"00", -- $0f7e8
          63465 => x"00", -- $0f7e9
          63466 => x"00", -- $0f7ea
          63467 => x"00", -- $0f7eb
          63468 => x"00", -- $0f7ec
          63469 => x"00", -- $0f7ed
          63470 => x"00", -- $0f7ee
          63471 => x"00", -- $0f7ef
          63472 => x"00", -- $0f7f0
          63473 => x"00", -- $0f7f1
          63474 => x"00", -- $0f7f2
          63475 => x"00", -- $0f7f3
          63476 => x"00", -- $0f7f4
          63477 => x"00", -- $0f7f5
          63478 => x"00", -- $0f7f6
          63479 => x"00", -- $0f7f7
          63480 => x"00", -- $0f7f8
          63481 => x"00", -- $0f7f9
          63482 => x"00", -- $0f7fa
          63483 => x"00", -- $0f7fb
          63484 => x"00", -- $0f7fc
          63485 => x"00", -- $0f7fd
          63486 => x"00", -- $0f7fe
          63487 => x"00", -- $0f7ff
          63488 => x"00", -- $0f800
          63489 => x"00", -- $0f801
          63490 => x"00", -- $0f802
          63491 => x"00", -- $0f803
          63492 => x"00", -- $0f804
          63493 => x"00", -- $0f805
          63494 => x"00", -- $0f806
          63495 => x"00", -- $0f807
          63496 => x"00", -- $0f808
          63497 => x"00", -- $0f809
          63498 => x"00", -- $0f80a
          63499 => x"00", -- $0f80b
          63500 => x"00", -- $0f80c
          63501 => x"00", -- $0f80d
          63502 => x"00", -- $0f80e
          63503 => x"00", -- $0f80f
          63504 => x"00", -- $0f810
          63505 => x"00", -- $0f811
          63506 => x"00", -- $0f812
          63507 => x"00", -- $0f813
          63508 => x"00", -- $0f814
          63509 => x"00", -- $0f815
          63510 => x"00", -- $0f816
          63511 => x"00", -- $0f817
          63512 => x"00", -- $0f818
          63513 => x"00", -- $0f819
          63514 => x"00", -- $0f81a
          63515 => x"00", -- $0f81b
          63516 => x"00", -- $0f81c
          63517 => x"00", -- $0f81d
          63518 => x"00", -- $0f81e
          63519 => x"00", -- $0f81f
          63520 => x"00", -- $0f820
          63521 => x"00", -- $0f821
          63522 => x"00", -- $0f822
          63523 => x"00", -- $0f823
          63524 => x"00", -- $0f824
          63525 => x"00", -- $0f825
          63526 => x"00", -- $0f826
          63527 => x"00", -- $0f827
          63528 => x"00", -- $0f828
          63529 => x"00", -- $0f829
          63530 => x"00", -- $0f82a
          63531 => x"00", -- $0f82b
          63532 => x"00", -- $0f82c
          63533 => x"00", -- $0f82d
          63534 => x"00", -- $0f82e
          63535 => x"00", -- $0f82f
          63536 => x"00", -- $0f830
          63537 => x"00", -- $0f831
          63538 => x"00", -- $0f832
          63539 => x"00", -- $0f833
          63540 => x"00", -- $0f834
          63541 => x"00", -- $0f835
          63542 => x"00", -- $0f836
          63543 => x"00", -- $0f837
          63544 => x"00", -- $0f838
          63545 => x"00", -- $0f839
          63546 => x"00", -- $0f83a
          63547 => x"00", -- $0f83b
          63548 => x"00", -- $0f83c
          63549 => x"00", -- $0f83d
          63550 => x"00", -- $0f83e
          63551 => x"00", -- $0f83f
          63552 => x"00", -- $0f840
          63553 => x"00", -- $0f841
          63554 => x"00", -- $0f842
          63555 => x"00", -- $0f843
          63556 => x"00", -- $0f844
          63557 => x"00", -- $0f845
          63558 => x"00", -- $0f846
          63559 => x"00", -- $0f847
          63560 => x"00", -- $0f848
          63561 => x"00", -- $0f849
          63562 => x"00", -- $0f84a
          63563 => x"00", -- $0f84b
          63564 => x"00", -- $0f84c
          63565 => x"00", -- $0f84d
          63566 => x"00", -- $0f84e
          63567 => x"00", -- $0f84f
          63568 => x"00", -- $0f850
          63569 => x"00", -- $0f851
          63570 => x"00", -- $0f852
          63571 => x"00", -- $0f853
          63572 => x"00", -- $0f854
          63573 => x"00", -- $0f855
          63574 => x"00", -- $0f856
          63575 => x"00", -- $0f857
          63576 => x"00", -- $0f858
          63577 => x"00", -- $0f859
          63578 => x"00", -- $0f85a
          63579 => x"00", -- $0f85b
          63580 => x"00", -- $0f85c
          63581 => x"00", -- $0f85d
          63582 => x"00", -- $0f85e
          63583 => x"00", -- $0f85f
          63584 => x"00", -- $0f860
          63585 => x"00", -- $0f861
          63586 => x"00", -- $0f862
          63587 => x"00", -- $0f863
          63588 => x"00", -- $0f864
          63589 => x"00", -- $0f865
          63590 => x"00", -- $0f866
          63591 => x"00", -- $0f867
          63592 => x"00", -- $0f868
          63593 => x"00", -- $0f869
          63594 => x"00", -- $0f86a
          63595 => x"00", -- $0f86b
          63596 => x"00", -- $0f86c
          63597 => x"00", -- $0f86d
          63598 => x"00", -- $0f86e
          63599 => x"00", -- $0f86f
          63600 => x"00", -- $0f870
          63601 => x"00", -- $0f871
          63602 => x"00", -- $0f872
          63603 => x"00", -- $0f873
          63604 => x"00", -- $0f874
          63605 => x"00", -- $0f875
          63606 => x"00", -- $0f876
          63607 => x"00", -- $0f877
          63608 => x"00", -- $0f878
          63609 => x"00", -- $0f879
          63610 => x"00", -- $0f87a
          63611 => x"00", -- $0f87b
          63612 => x"00", -- $0f87c
          63613 => x"00", -- $0f87d
          63614 => x"00", -- $0f87e
          63615 => x"00", -- $0f87f
          63616 => x"00", -- $0f880
          63617 => x"00", -- $0f881
          63618 => x"00", -- $0f882
          63619 => x"00", -- $0f883
          63620 => x"00", -- $0f884
          63621 => x"00", -- $0f885
          63622 => x"00", -- $0f886
          63623 => x"00", -- $0f887
          63624 => x"00", -- $0f888
          63625 => x"00", -- $0f889
          63626 => x"00", -- $0f88a
          63627 => x"00", -- $0f88b
          63628 => x"00", -- $0f88c
          63629 => x"00", -- $0f88d
          63630 => x"00", -- $0f88e
          63631 => x"00", -- $0f88f
          63632 => x"00", -- $0f890
          63633 => x"00", -- $0f891
          63634 => x"00", -- $0f892
          63635 => x"00", -- $0f893
          63636 => x"00", -- $0f894
          63637 => x"00", -- $0f895
          63638 => x"00", -- $0f896
          63639 => x"00", -- $0f897
          63640 => x"00", -- $0f898
          63641 => x"00", -- $0f899
          63642 => x"00", -- $0f89a
          63643 => x"00", -- $0f89b
          63644 => x"00", -- $0f89c
          63645 => x"00", -- $0f89d
          63646 => x"00", -- $0f89e
          63647 => x"00", -- $0f89f
          63648 => x"00", -- $0f8a0
          63649 => x"00", -- $0f8a1
          63650 => x"00", -- $0f8a2
          63651 => x"00", -- $0f8a3
          63652 => x"00", -- $0f8a4
          63653 => x"00", -- $0f8a5
          63654 => x"00", -- $0f8a6
          63655 => x"00", -- $0f8a7
          63656 => x"00", -- $0f8a8
          63657 => x"00", -- $0f8a9
          63658 => x"00", -- $0f8aa
          63659 => x"00", -- $0f8ab
          63660 => x"00", -- $0f8ac
          63661 => x"00", -- $0f8ad
          63662 => x"00", -- $0f8ae
          63663 => x"00", -- $0f8af
          63664 => x"00", -- $0f8b0
          63665 => x"00", -- $0f8b1
          63666 => x"00", -- $0f8b2
          63667 => x"00", -- $0f8b3
          63668 => x"00", -- $0f8b4
          63669 => x"00", -- $0f8b5
          63670 => x"00", -- $0f8b6
          63671 => x"00", -- $0f8b7
          63672 => x"00", -- $0f8b8
          63673 => x"00", -- $0f8b9
          63674 => x"00", -- $0f8ba
          63675 => x"00", -- $0f8bb
          63676 => x"00", -- $0f8bc
          63677 => x"00", -- $0f8bd
          63678 => x"00", -- $0f8be
          63679 => x"00", -- $0f8bf
          63680 => x"00", -- $0f8c0
          63681 => x"00", -- $0f8c1
          63682 => x"00", -- $0f8c2
          63683 => x"00", -- $0f8c3
          63684 => x"00", -- $0f8c4
          63685 => x"00", -- $0f8c5
          63686 => x"00", -- $0f8c6
          63687 => x"00", -- $0f8c7
          63688 => x"00", -- $0f8c8
          63689 => x"00", -- $0f8c9
          63690 => x"00", -- $0f8ca
          63691 => x"00", -- $0f8cb
          63692 => x"00", -- $0f8cc
          63693 => x"00", -- $0f8cd
          63694 => x"00", -- $0f8ce
          63695 => x"00", -- $0f8cf
          63696 => x"00", -- $0f8d0
          63697 => x"00", -- $0f8d1
          63698 => x"00", -- $0f8d2
          63699 => x"00", -- $0f8d3
          63700 => x"00", -- $0f8d4
          63701 => x"00", -- $0f8d5
          63702 => x"00", -- $0f8d6
          63703 => x"00", -- $0f8d7
          63704 => x"00", -- $0f8d8
          63705 => x"00", -- $0f8d9
          63706 => x"00", -- $0f8da
          63707 => x"00", -- $0f8db
          63708 => x"00", -- $0f8dc
          63709 => x"00", -- $0f8dd
          63710 => x"00", -- $0f8de
          63711 => x"00", -- $0f8df
          63712 => x"00", -- $0f8e0
          63713 => x"00", -- $0f8e1
          63714 => x"00", -- $0f8e2
          63715 => x"00", -- $0f8e3
          63716 => x"00", -- $0f8e4
          63717 => x"00", -- $0f8e5
          63718 => x"00", -- $0f8e6
          63719 => x"00", -- $0f8e7
          63720 => x"00", -- $0f8e8
          63721 => x"00", -- $0f8e9
          63722 => x"00", -- $0f8ea
          63723 => x"00", -- $0f8eb
          63724 => x"00", -- $0f8ec
          63725 => x"00", -- $0f8ed
          63726 => x"00", -- $0f8ee
          63727 => x"00", -- $0f8ef
          63728 => x"00", -- $0f8f0
          63729 => x"00", -- $0f8f1
          63730 => x"00", -- $0f8f2
          63731 => x"00", -- $0f8f3
          63732 => x"00", -- $0f8f4
          63733 => x"00", -- $0f8f5
          63734 => x"00", -- $0f8f6
          63735 => x"00", -- $0f8f7
          63736 => x"00", -- $0f8f8
          63737 => x"00", -- $0f8f9
          63738 => x"00", -- $0f8fa
          63739 => x"00", -- $0f8fb
          63740 => x"00", -- $0f8fc
          63741 => x"00", -- $0f8fd
          63742 => x"00", -- $0f8fe
          63743 => x"00", -- $0f8ff
          63744 => x"00", -- $0f900
          63745 => x"00", -- $0f901
          63746 => x"00", -- $0f902
          63747 => x"00", -- $0f903
          63748 => x"00", -- $0f904
          63749 => x"00", -- $0f905
          63750 => x"00", -- $0f906
          63751 => x"00", -- $0f907
          63752 => x"00", -- $0f908
          63753 => x"00", -- $0f909
          63754 => x"00", -- $0f90a
          63755 => x"00", -- $0f90b
          63756 => x"00", -- $0f90c
          63757 => x"00", -- $0f90d
          63758 => x"00", -- $0f90e
          63759 => x"00", -- $0f90f
          63760 => x"00", -- $0f910
          63761 => x"00", -- $0f911
          63762 => x"00", -- $0f912
          63763 => x"00", -- $0f913
          63764 => x"00", -- $0f914
          63765 => x"00", -- $0f915
          63766 => x"00", -- $0f916
          63767 => x"00", -- $0f917
          63768 => x"00", -- $0f918
          63769 => x"00", -- $0f919
          63770 => x"00", -- $0f91a
          63771 => x"00", -- $0f91b
          63772 => x"00", -- $0f91c
          63773 => x"00", -- $0f91d
          63774 => x"00", -- $0f91e
          63775 => x"00", -- $0f91f
          63776 => x"00", -- $0f920
          63777 => x"00", -- $0f921
          63778 => x"00", -- $0f922
          63779 => x"00", -- $0f923
          63780 => x"00", -- $0f924
          63781 => x"00", -- $0f925
          63782 => x"00", -- $0f926
          63783 => x"00", -- $0f927
          63784 => x"00", -- $0f928
          63785 => x"00", -- $0f929
          63786 => x"00", -- $0f92a
          63787 => x"00", -- $0f92b
          63788 => x"00", -- $0f92c
          63789 => x"00", -- $0f92d
          63790 => x"00", -- $0f92e
          63791 => x"00", -- $0f92f
          63792 => x"00", -- $0f930
          63793 => x"00", -- $0f931
          63794 => x"00", -- $0f932
          63795 => x"00", -- $0f933
          63796 => x"00", -- $0f934
          63797 => x"00", -- $0f935
          63798 => x"00", -- $0f936
          63799 => x"00", -- $0f937
          63800 => x"00", -- $0f938
          63801 => x"00", -- $0f939
          63802 => x"00", -- $0f93a
          63803 => x"00", -- $0f93b
          63804 => x"00", -- $0f93c
          63805 => x"00", -- $0f93d
          63806 => x"00", -- $0f93e
          63807 => x"00", -- $0f93f
          63808 => x"00", -- $0f940
          63809 => x"00", -- $0f941
          63810 => x"00", -- $0f942
          63811 => x"00", -- $0f943
          63812 => x"00", -- $0f944
          63813 => x"00", -- $0f945
          63814 => x"00", -- $0f946
          63815 => x"00", -- $0f947
          63816 => x"00", -- $0f948
          63817 => x"00", -- $0f949
          63818 => x"00", -- $0f94a
          63819 => x"00", -- $0f94b
          63820 => x"00", -- $0f94c
          63821 => x"00", -- $0f94d
          63822 => x"00", -- $0f94e
          63823 => x"00", -- $0f94f
          63824 => x"00", -- $0f950
          63825 => x"00", -- $0f951
          63826 => x"00", -- $0f952
          63827 => x"00", -- $0f953
          63828 => x"00", -- $0f954
          63829 => x"00", -- $0f955
          63830 => x"00", -- $0f956
          63831 => x"00", -- $0f957
          63832 => x"00", -- $0f958
          63833 => x"00", -- $0f959
          63834 => x"00", -- $0f95a
          63835 => x"00", -- $0f95b
          63836 => x"00", -- $0f95c
          63837 => x"00", -- $0f95d
          63838 => x"00", -- $0f95e
          63839 => x"00", -- $0f95f
          63840 => x"00", -- $0f960
          63841 => x"00", -- $0f961
          63842 => x"00", -- $0f962
          63843 => x"00", -- $0f963
          63844 => x"00", -- $0f964
          63845 => x"00", -- $0f965
          63846 => x"00", -- $0f966
          63847 => x"00", -- $0f967
          63848 => x"00", -- $0f968
          63849 => x"00", -- $0f969
          63850 => x"00", -- $0f96a
          63851 => x"00", -- $0f96b
          63852 => x"00", -- $0f96c
          63853 => x"00", -- $0f96d
          63854 => x"00", -- $0f96e
          63855 => x"00", -- $0f96f
          63856 => x"00", -- $0f970
          63857 => x"00", -- $0f971
          63858 => x"00", -- $0f972
          63859 => x"00", -- $0f973
          63860 => x"00", -- $0f974
          63861 => x"00", -- $0f975
          63862 => x"00", -- $0f976
          63863 => x"00", -- $0f977
          63864 => x"00", -- $0f978
          63865 => x"00", -- $0f979
          63866 => x"00", -- $0f97a
          63867 => x"00", -- $0f97b
          63868 => x"00", -- $0f97c
          63869 => x"00", -- $0f97d
          63870 => x"00", -- $0f97e
          63871 => x"00", -- $0f97f
          63872 => x"00", -- $0f980
          63873 => x"00", -- $0f981
          63874 => x"00", -- $0f982
          63875 => x"00", -- $0f983
          63876 => x"00", -- $0f984
          63877 => x"00", -- $0f985
          63878 => x"00", -- $0f986
          63879 => x"00", -- $0f987
          63880 => x"00", -- $0f988
          63881 => x"00", -- $0f989
          63882 => x"00", -- $0f98a
          63883 => x"00", -- $0f98b
          63884 => x"00", -- $0f98c
          63885 => x"00", -- $0f98d
          63886 => x"00", -- $0f98e
          63887 => x"00", -- $0f98f
          63888 => x"00", -- $0f990
          63889 => x"00", -- $0f991
          63890 => x"00", -- $0f992
          63891 => x"00", -- $0f993
          63892 => x"00", -- $0f994
          63893 => x"00", -- $0f995
          63894 => x"00", -- $0f996
          63895 => x"00", -- $0f997
          63896 => x"00", -- $0f998
          63897 => x"00", -- $0f999
          63898 => x"00", -- $0f99a
          63899 => x"00", -- $0f99b
          63900 => x"00", -- $0f99c
          63901 => x"00", -- $0f99d
          63902 => x"00", -- $0f99e
          63903 => x"00", -- $0f99f
          63904 => x"00", -- $0f9a0
          63905 => x"00", -- $0f9a1
          63906 => x"00", -- $0f9a2
          63907 => x"00", -- $0f9a3
          63908 => x"00", -- $0f9a4
          63909 => x"00", -- $0f9a5
          63910 => x"00", -- $0f9a6
          63911 => x"00", -- $0f9a7
          63912 => x"00", -- $0f9a8
          63913 => x"00", -- $0f9a9
          63914 => x"00", -- $0f9aa
          63915 => x"00", -- $0f9ab
          63916 => x"00", -- $0f9ac
          63917 => x"00", -- $0f9ad
          63918 => x"00", -- $0f9ae
          63919 => x"00", -- $0f9af
          63920 => x"00", -- $0f9b0
          63921 => x"00", -- $0f9b1
          63922 => x"00", -- $0f9b2
          63923 => x"00", -- $0f9b3
          63924 => x"00", -- $0f9b4
          63925 => x"00", -- $0f9b5
          63926 => x"00", -- $0f9b6
          63927 => x"00", -- $0f9b7
          63928 => x"00", -- $0f9b8
          63929 => x"00", -- $0f9b9
          63930 => x"00", -- $0f9ba
          63931 => x"00", -- $0f9bb
          63932 => x"00", -- $0f9bc
          63933 => x"00", -- $0f9bd
          63934 => x"00", -- $0f9be
          63935 => x"00", -- $0f9bf
          63936 => x"00", -- $0f9c0
          63937 => x"00", -- $0f9c1
          63938 => x"00", -- $0f9c2
          63939 => x"00", -- $0f9c3
          63940 => x"00", -- $0f9c4
          63941 => x"00", -- $0f9c5
          63942 => x"00", -- $0f9c6
          63943 => x"00", -- $0f9c7
          63944 => x"00", -- $0f9c8
          63945 => x"00", -- $0f9c9
          63946 => x"00", -- $0f9ca
          63947 => x"00", -- $0f9cb
          63948 => x"00", -- $0f9cc
          63949 => x"00", -- $0f9cd
          63950 => x"00", -- $0f9ce
          63951 => x"00", -- $0f9cf
          63952 => x"00", -- $0f9d0
          63953 => x"00", -- $0f9d1
          63954 => x"00", -- $0f9d2
          63955 => x"00", -- $0f9d3
          63956 => x"00", -- $0f9d4
          63957 => x"00", -- $0f9d5
          63958 => x"00", -- $0f9d6
          63959 => x"00", -- $0f9d7
          63960 => x"00", -- $0f9d8
          63961 => x"00", -- $0f9d9
          63962 => x"00", -- $0f9da
          63963 => x"00", -- $0f9db
          63964 => x"00", -- $0f9dc
          63965 => x"00", -- $0f9dd
          63966 => x"00", -- $0f9de
          63967 => x"00", -- $0f9df
          63968 => x"00", -- $0f9e0
          63969 => x"00", -- $0f9e1
          63970 => x"00", -- $0f9e2
          63971 => x"00", -- $0f9e3
          63972 => x"00", -- $0f9e4
          63973 => x"00", -- $0f9e5
          63974 => x"00", -- $0f9e6
          63975 => x"00", -- $0f9e7
          63976 => x"00", -- $0f9e8
          63977 => x"00", -- $0f9e9
          63978 => x"00", -- $0f9ea
          63979 => x"00", -- $0f9eb
          63980 => x"00", -- $0f9ec
          63981 => x"00", -- $0f9ed
          63982 => x"00", -- $0f9ee
          63983 => x"00", -- $0f9ef
          63984 => x"00", -- $0f9f0
          63985 => x"00", -- $0f9f1
          63986 => x"00", -- $0f9f2
          63987 => x"00", -- $0f9f3
          63988 => x"00", -- $0f9f4
          63989 => x"00", -- $0f9f5
          63990 => x"00", -- $0f9f6
          63991 => x"00", -- $0f9f7
          63992 => x"00", -- $0f9f8
          63993 => x"00", -- $0f9f9
          63994 => x"00", -- $0f9fa
          63995 => x"00", -- $0f9fb
          63996 => x"00", -- $0f9fc
          63997 => x"00", -- $0f9fd
          63998 => x"00", -- $0f9fe
          63999 => x"00", -- $0f9ff
          64000 => x"00", -- $0fa00
          64001 => x"00", -- $0fa01
          64002 => x"00", -- $0fa02
          64003 => x"00", -- $0fa03
          64004 => x"00", -- $0fa04
          64005 => x"00", -- $0fa05
          64006 => x"00", -- $0fa06
          64007 => x"00", -- $0fa07
          64008 => x"00", -- $0fa08
          64009 => x"00", -- $0fa09
          64010 => x"00", -- $0fa0a
          64011 => x"00", -- $0fa0b
          64012 => x"00", -- $0fa0c
          64013 => x"00", -- $0fa0d
          64014 => x"00", -- $0fa0e
          64015 => x"00", -- $0fa0f
          64016 => x"00", -- $0fa10
          64017 => x"00", -- $0fa11
          64018 => x"00", -- $0fa12
          64019 => x"00", -- $0fa13
          64020 => x"00", -- $0fa14
          64021 => x"00", -- $0fa15
          64022 => x"00", -- $0fa16
          64023 => x"00", -- $0fa17
          64024 => x"00", -- $0fa18
          64025 => x"00", -- $0fa19
          64026 => x"00", -- $0fa1a
          64027 => x"00", -- $0fa1b
          64028 => x"00", -- $0fa1c
          64029 => x"00", -- $0fa1d
          64030 => x"00", -- $0fa1e
          64031 => x"00", -- $0fa1f
          64032 => x"00", -- $0fa20
          64033 => x"00", -- $0fa21
          64034 => x"00", -- $0fa22
          64035 => x"00", -- $0fa23
          64036 => x"00", -- $0fa24
          64037 => x"00", -- $0fa25
          64038 => x"00", -- $0fa26
          64039 => x"00", -- $0fa27
          64040 => x"00", -- $0fa28
          64041 => x"00", -- $0fa29
          64042 => x"00", -- $0fa2a
          64043 => x"00", -- $0fa2b
          64044 => x"00", -- $0fa2c
          64045 => x"00", -- $0fa2d
          64046 => x"00", -- $0fa2e
          64047 => x"00", -- $0fa2f
          64048 => x"00", -- $0fa30
          64049 => x"00", -- $0fa31
          64050 => x"00", -- $0fa32
          64051 => x"00", -- $0fa33
          64052 => x"00", -- $0fa34
          64053 => x"00", -- $0fa35
          64054 => x"00", -- $0fa36
          64055 => x"00", -- $0fa37
          64056 => x"00", -- $0fa38
          64057 => x"00", -- $0fa39
          64058 => x"00", -- $0fa3a
          64059 => x"00", -- $0fa3b
          64060 => x"00", -- $0fa3c
          64061 => x"00", -- $0fa3d
          64062 => x"00", -- $0fa3e
          64063 => x"00", -- $0fa3f
          64064 => x"00", -- $0fa40
          64065 => x"00", -- $0fa41
          64066 => x"00", -- $0fa42
          64067 => x"00", -- $0fa43
          64068 => x"00", -- $0fa44
          64069 => x"00", -- $0fa45
          64070 => x"00", -- $0fa46
          64071 => x"00", -- $0fa47
          64072 => x"00", -- $0fa48
          64073 => x"00", -- $0fa49
          64074 => x"00", -- $0fa4a
          64075 => x"00", -- $0fa4b
          64076 => x"00", -- $0fa4c
          64077 => x"00", -- $0fa4d
          64078 => x"00", -- $0fa4e
          64079 => x"00", -- $0fa4f
          64080 => x"00", -- $0fa50
          64081 => x"00", -- $0fa51
          64082 => x"00", -- $0fa52
          64083 => x"00", -- $0fa53
          64084 => x"00", -- $0fa54
          64085 => x"00", -- $0fa55
          64086 => x"00", -- $0fa56
          64087 => x"00", -- $0fa57
          64088 => x"00", -- $0fa58
          64089 => x"00", -- $0fa59
          64090 => x"00", -- $0fa5a
          64091 => x"00", -- $0fa5b
          64092 => x"00", -- $0fa5c
          64093 => x"00", -- $0fa5d
          64094 => x"00", -- $0fa5e
          64095 => x"00", -- $0fa5f
          64096 => x"00", -- $0fa60
          64097 => x"00", -- $0fa61
          64098 => x"00", -- $0fa62
          64099 => x"00", -- $0fa63
          64100 => x"00", -- $0fa64
          64101 => x"00", -- $0fa65
          64102 => x"00", -- $0fa66
          64103 => x"00", -- $0fa67
          64104 => x"00", -- $0fa68
          64105 => x"00", -- $0fa69
          64106 => x"00", -- $0fa6a
          64107 => x"00", -- $0fa6b
          64108 => x"00", -- $0fa6c
          64109 => x"00", -- $0fa6d
          64110 => x"00", -- $0fa6e
          64111 => x"00", -- $0fa6f
          64112 => x"00", -- $0fa70
          64113 => x"00", -- $0fa71
          64114 => x"00", -- $0fa72
          64115 => x"00", -- $0fa73
          64116 => x"00", -- $0fa74
          64117 => x"00", -- $0fa75
          64118 => x"00", -- $0fa76
          64119 => x"00", -- $0fa77
          64120 => x"00", -- $0fa78
          64121 => x"00", -- $0fa79
          64122 => x"00", -- $0fa7a
          64123 => x"00", -- $0fa7b
          64124 => x"00", -- $0fa7c
          64125 => x"00", -- $0fa7d
          64126 => x"00", -- $0fa7e
          64127 => x"00", -- $0fa7f
          64128 => x"00", -- $0fa80
          64129 => x"00", -- $0fa81
          64130 => x"00", -- $0fa82
          64131 => x"00", -- $0fa83
          64132 => x"00", -- $0fa84
          64133 => x"00", -- $0fa85
          64134 => x"00", -- $0fa86
          64135 => x"00", -- $0fa87
          64136 => x"00", -- $0fa88
          64137 => x"00", -- $0fa89
          64138 => x"00", -- $0fa8a
          64139 => x"00", -- $0fa8b
          64140 => x"00", -- $0fa8c
          64141 => x"00", -- $0fa8d
          64142 => x"00", -- $0fa8e
          64143 => x"00", -- $0fa8f
          64144 => x"00", -- $0fa90
          64145 => x"00", -- $0fa91
          64146 => x"00", -- $0fa92
          64147 => x"00", -- $0fa93
          64148 => x"00", -- $0fa94
          64149 => x"00", -- $0fa95
          64150 => x"00", -- $0fa96
          64151 => x"00", -- $0fa97
          64152 => x"00", -- $0fa98
          64153 => x"00", -- $0fa99
          64154 => x"00", -- $0fa9a
          64155 => x"00", -- $0fa9b
          64156 => x"00", -- $0fa9c
          64157 => x"00", -- $0fa9d
          64158 => x"00", -- $0fa9e
          64159 => x"00", -- $0fa9f
          64160 => x"00", -- $0faa0
          64161 => x"00", -- $0faa1
          64162 => x"00", -- $0faa2
          64163 => x"00", -- $0faa3
          64164 => x"00", -- $0faa4
          64165 => x"00", -- $0faa5
          64166 => x"00", -- $0faa6
          64167 => x"00", -- $0faa7
          64168 => x"00", -- $0faa8
          64169 => x"00", -- $0faa9
          64170 => x"00", -- $0faaa
          64171 => x"00", -- $0faab
          64172 => x"00", -- $0faac
          64173 => x"00", -- $0faad
          64174 => x"00", -- $0faae
          64175 => x"00", -- $0faaf
          64176 => x"00", -- $0fab0
          64177 => x"00", -- $0fab1
          64178 => x"00", -- $0fab2
          64179 => x"00", -- $0fab3
          64180 => x"00", -- $0fab4
          64181 => x"00", -- $0fab5
          64182 => x"00", -- $0fab6
          64183 => x"00", -- $0fab7
          64184 => x"00", -- $0fab8
          64185 => x"00", -- $0fab9
          64186 => x"00", -- $0faba
          64187 => x"00", -- $0fabb
          64188 => x"00", -- $0fabc
          64189 => x"00", -- $0fabd
          64190 => x"00", -- $0fabe
          64191 => x"00", -- $0fabf
          64192 => x"00", -- $0fac0
          64193 => x"00", -- $0fac1
          64194 => x"00", -- $0fac2
          64195 => x"00", -- $0fac3
          64196 => x"00", -- $0fac4
          64197 => x"00", -- $0fac5
          64198 => x"00", -- $0fac6
          64199 => x"00", -- $0fac7
          64200 => x"00", -- $0fac8
          64201 => x"00", -- $0fac9
          64202 => x"00", -- $0faca
          64203 => x"00", -- $0facb
          64204 => x"00", -- $0facc
          64205 => x"00", -- $0facd
          64206 => x"00", -- $0face
          64207 => x"00", -- $0facf
          64208 => x"00", -- $0fad0
          64209 => x"00", -- $0fad1
          64210 => x"00", -- $0fad2
          64211 => x"00", -- $0fad3
          64212 => x"00", -- $0fad4
          64213 => x"00", -- $0fad5
          64214 => x"00", -- $0fad6
          64215 => x"00", -- $0fad7
          64216 => x"00", -- $0fad8
          64217 => x"00", -- $0fad9
          64218 => x"00", -- $0fada
          64219 => x"00", -- $0fadb
          64220 => x"00", -- $0fadc
          64221 => x"00", -- $0fadd
          64222 => x"00", -- $0fade
          64223 => x"00", -- $0fadf
          64224 => x"00", -- $0fae0
          64225 => x"00", -- $0fae1
          64226 => x"00", -- $0fae2
          64227 => x"00", -- $0fae3
          64228 => x"00", -- $0fae4
          64229 => x"00", -- $0fae5
          64230 => x"00", -- $0fae6
          64231 => x"00", -- $0fae7
          64232 => x"00", -- $0fae8
          64233 => x"00", -- $0fae9
          64234 => x"00", -- $0faea
          64235 => x"00", -- $0faeb
          64236 => x"00", -- $0faec
          64237 => x"00", -- $0faed
          64238 => x"00", -- $0faee
          64239 => x"00", -- $0faef
          64240 => x"00", -- $0faf0
          64241 => x"00", -- $0faf1
          64242 => x"00", -- $0faf2
          64243 => x"00", -- $0faf3
          64244 => x"00", -- $0faf4
          64245 => x"00", -- $0faf5
          64246 => x"00", -- $0faf6
          64247 => x"00", -- $0faf7
          64248 => x"00", -- $0faf8
          64249 => x"00", -- $0faf9
          64250 => x"00", -- $0fafa
          64251 => x"00", -- $0fafb
          64252 => x"00", -- $0fafc
          64253 => x"00", -- $0fafd
          64254 => x"00", -- $0fafe
          64255 => x"00", -- $0faff
          64256 => x"00", -- $0fb00
          64257 => x"00", -- $0fb01
          64258 => x"00", -- $0fb02
          64259 => x"00", -- $0fb03
          64260 => x"00", -- $0fb04
          64261 => x"00", -- $0fb05
          64262 => x"00", -- $0fb06
          64263 => x"00", -- $0fb07
          64264 => x"00", -- $0fb08
          64265 => x"00", -- $0fb09
          64266 => x"00", -- $0fb0a
          64267 => x"00", -- $0fb0b
          64268 => x"00", -- $0fb0c
          64269 => x"00", -- $0fb0d
          64270 => x"00", -- $0fb0e
          64271 => x"00", -- $0fb0f
          64272 => x"00", -- $0fb10
          64273 => x"00", -- $0fb11
          64274 => x"00", -- $0fb12
          64275 => x"00", -- $0fb13
          64276 => x"00", -- $0fb14
          64277 => x"00", -- $0fb15
          64278 => x"00", -- $0fb16
          64279 => x"00", -- $0fb17
          64280 => x"00", -- $0fb18
          64281 => x"00", -- $0fb19
          64282 => x"00", -- $0fb1a
          64283 => x"00", -- $0fb1b
          64284 => x"00", -- $0fb1c
          64285 => x"00", -- $0fb1d
          64286 => x"00", -- $0fb1e
          64287 => x"00", -- $0fb1f
          64288 => x"00", -- $0fb20
          64289 => x"00", -- $0fb21
          64290 => x"00", -- $0fb22
          64291 => x"00", -- $0fb23
          64292 => x"00", -- $0fb24
          64293 => x"00", -- $0fb25
          64294 => x"00", -- $0fb26
          64295 => x"00", -- $0fb27
          64296 => x"00", -- $0fb28
          64297 => x"00", -- $0fb29
          64298 => x"00", -- $0fb2a
          64299 => x"00", -- $0fb2b
          64300 => x"00", -- $0fb2c
          64301 => x"00", -- $0fb2d
          64302 => x"00", -- $0fb2e
          64303 => x"00", -- $0fb2f
          64304 => x"00", -- $0fb30
          64305 => x"00", -- $0fb31
          64306 => x"00", -- $0fb32
          64307 => x"00", -- $0fb33
          64308 => x"00", -- $0fb34
          64309 => x"00", -- $0fb35
          64310 => x"00", -- $0fb36
          64311 => x"00", -- $0fb37
          64312 => x"00", -- $0fb38
          64313 => x"00", -- $0fb39
          64314 => x"00", -- $0fb3a
          64315 => x"00", -- $0fb3b
          64316 => x"00", -- $0fb3c
          64317 => x"00", -- $0fb3d
          64318 => x"00", -- $0fb3e
          64319 => x"00", -- $0fb3f
          64320 => x"00", -- $0fb40
          64321 => x"00", -- $0fb41
          64322 => x"00", -- $0fb42
          64323 => x"00", -- $0fb43
          64324 => x"00", -- $0fb44
          64325 => x"00", -- $0fb45
          64326 => x"00", -- $0fb46
          64327 => x"00", -- $0fb47
          64328 => x"00", -- $0fb48
          64329 => x"00", -- $0fb49
          64330 => x"00", -- $0fb4a
          64331 => x"00", -- $0fb4b
          64332 => x"00", -- $0fb4c
          64333 => x"00", -- $0fb4d
          64334 => x"00", -- $0fb4e
          64335 => x"00", -- $0fb4f
          64336 => x"00", -- $0fb50
          64337 => x"00", -- $0fb51
          64338 => x"00", -- $0fb52
          64339 => x"00", -- $0fb53
          64340 => x"00", -- $0fb54
          64341 => x"00", -- $0fb55
          64342 => x"00", -- $0fb56
          64343 => x"00", -- $0fb57
          64344 => x"00", -- $0fb58
          64345 => x"00", -- $0fb59
          64346 => x"00", -- $0fb5a
          64347 => x"00", -- $0fb5b
          64348 => x"00", -- $0fb5c
          64349 => x"00", -- $0fb5d
          64350 => x"00", -- $0fb5e
          64351 => x"00", -- $0fb5f
          64352 => x"00", -- $0fb60
          64353 => x"00", -- $0fb61
          64354 => x"00", -- $0fb62
          64355 => x"00", -- $0fb63
          64356 => x"00", -- $0fb64
          64357 => x"00", -- $0fb65
          64358 => x"00", -- $0fb66
          64359 => x"00", -- $0fb67
          64360 => x"00", -- $0fb68
          64361 => x"00", -- $0fb69
          64362 => x"00", -- $0fb6a
          64363 => x"00", -- $0fb6b
          64364 => x"00", -- $0fb6c
          64365 => x"00", -- $0fb6d
          64366 => x"00", -- $0fb6e
          64367 => x"00", -- $0fb6f
          64368 => x"00", -- $0fb70
          64369 => x"00", -- $0fb71
          64370 => x"00", -- $0fb72
          64371 => x"00", -- $0fb73
          64372 => x"00", -- $0fb74
          64373 => x"00", -- $0fb75
          64374 => x"00", -- $0fb76
          64375 => x"00", -- $0fb77
          64376 => x"00", -- $0fb78
          64377 => x"00", -- $0fb79
          64378 => x"00", -- $0fb7a
          64379 => x"00", -- $0fb7b
          64380 => x"00", -- $0fb7c
          64381 => x"00", -- $0fb7d
          64382 => x"00", -- $0fb7e
          64383 => x"00", -- $0fb7f
          64384 => x"00", -- $0fb80
          64385 => x"00", -- $0fb81
          64386 => x"00", -- $0fb82
          64387 => x"00", -- $0fb83
          64388 => x"00", -- $0fb84
          64389 => x"00", -- $0fb85
          64390 => x"00", -- $0fb86
          64391 => x"00", -- $0fb87
          64392 => x"00", -- $0fb88
          64393 => x"00", -- $0fb89
          64394 => x"00", -- $0fb8a
          64395 => x"00", -- $0fb8b
          64396 => x"00", -- $0fb8c
          64397 => x"00", -- $0fb8d
          64398 => x"00", -- $0fb8e
          64399 => x"00", -- $0fb8f
          64400 => x"00", -- $0fb90
          64401 => x"00", -- $0fb91
          64402 => x"00", -- $0fb92
          64403 => x"00", -- $0fb93
          64404 => x"00", -- $0fb94
          64405 => x"00", -- $0fb95
          64406 => x"00", -- $0fb96
          64407 => x"00", -- $0fb97
          64408 => x"00", -- $0fb98
          64409 => x"00", -- $0fb99
          64410 => x"00", -- $0fb9a
          64411 => x"00", -- $0fb9b
          64412 => x"00", -- $0fb9c
          64413 => x"00", -- $0fb9d
          64414 => x"00", -- $0fb9e
          64415 => x"00", -- $0fb9f
          64416 => x"00", -- $0fba0
          64417 => x"00", -- $0fba1
          64418 => x"00", -- $0fba2
          64419 => x"00", -- $0fba3
          64420 => x"00", -- $0fba4
          64421 => x"00", -- $0fba5
          64422 => x"00", -- $0fba6
          64423 => x"00", -- $0fba7
          64424 => x"00", -- $0fba8
          64425 => x"00", -- $0fba9
          64426 => x"00", -- $0fbaa
          64427 => x"00", -- $0fbab
          64428 => x"00", -- $0fbac
          64429 => x"00", -- $0fbad
          64430 => x"00", -- $0fbae
          64431 => x"00", -- $0fbaf
          64432 => x"00", -- $0fbb0
          64433 => x"00", -- $0fbb1
          64434 => x"00", -- $0fbb2
          64435 => x"00", -- $0fbb3
          64436 => x"00", -- $0fbb4
          64437 => x"00", -- $0fbb5
          64438 => x"00", -- $0fbb6
          64439 => x"00", -- $0fbb7
          64440 => x"00", -- $0fbb8
          64441 => x"00", -- $0fbb9
          64442 => x"00", -- $0fbba
          64443 => x"00", -- $0fbbb
          64444 => x"00", -- $0fbbc
          64445 => x"00", -- $0fbbd
          64446 => x"00", -- $0fbbe
          64447 => x"00", -- $0fbbf
          64448 => x"00", -- $0fbc0
          64449 => x"00", -- $0fbc1
          64450 => x"00", -- $0fbc2
          64451 => x"00", -- $0fbc3
          64452 => x"00", -- $0fbc4
          64453 => x"00", -- $0fbc5
          64454 => x"00", -- $0fbc6
          64455 => x"00", -- $0fbc7
          64456 => x"00", -- $0fbc8
          64457 => x"00", -- $0fbc9
          64458 => x"00", -- $0fbca
          64459 => x"00", -- $0fbcb
          64460 => x"00", -- $0fbcc
          64461 => x"00", -- $0fbcd
          64462 => x"00", -- $0fbce
          64463 => x"00", -- $0fbcf
          64464 => x"00", -- $0fbd0
          64465 => x"00", -- $0fbd1
          64466 => x"00", -- $0fbd2
          64467 => x"00", -- $0fbd3
          64468 => x"00", -- $0fbd4
          64469 => x"00", -- $0fbd5
          64470 => x"00", -- $0fbd6
          64471 => x"00", -- $0fbd7
          64472 => x"00", -- $0fbd8
          64473 => x"00", -- $0fbd9
          64474 => x"00", -- $0fbda
          64475 => x"00", -- $0fbdb
          64476 => x"00", -- $0fbdc
          64477 => x"00", -- $0fbdd
          64478 => x"00", -- $0fbde
          64479 => x"00", -- $0fbdf
          64480 => x"00", -- $0fbe0
          64481 => x"00", -- $0fbe1
          64482 => x"00", -- $0fbe2
          64483 => x"00", -- $0fbe3
          64484 => x"00", -- $0fbe4
          64485 => x"00", -- $0fbe5
          64486 => x"00", -- $0fbe6
          64487 => x"00", -- $0fbe7
          64488 => x"00", -- $0fbe8
          64489 => x"00", -- $0fbe9
          64490 => x"00", -- $0fbea
          64491 => x"00", -- $0fbeb
          64492 => x"00", -- $0fbec
          64493 => x"00", -- $0fbed
          64494 => x"00", -- $0fbee
          64495 => x"00", -- $0fbef
          64496 => x"00", -- $0fbf0
          64497 => x"00", -- $0fbf1
          64498 => x"00", -- $0fbf2
          64499 => x"00", -- $0fbf3
          64500 => x"00", -- $0fbf4
          64501 => x"00", -- $0fbf5
          64502 => x"00", -- $0fbf6
          64503 => x"00", -- $0fbf7
          64504 => x"00", -- $0fbf8
          64505 => x"00", -- $0fbf9
          64506 => x"00", -- $0fbfa
          64507 => x"00", -- $0fbfb
          64508 => x"00", -- $0fbfc
          64509 => x"00", -- $0fbfd
          64510 => x"00", -- $0fbfe
          64511 => x"00", -- $0fbff
          64512 => x"00", -- $0fc00
          64513 => x"00", -- $0fc01
          64514 => x"00", -- $0fc02
          64515 => x"00", -- $0fc03
          64516 => x"00", -- $0fc04
          64517 => x"00", -- $0fc05
          64518 => x"00", -- $0fc06
          64519 => x"00", -- $0fc07
          64520 => x"00", -- $0fc08
          64521 => x"00", -- $0fc09
          64522 => x"00", -- $0fc0a
          64523 => x"00", -- $0fc0b
          64524 => x"00", -- $0fc0c
          64525 => x"00", -- $0fc0d
          64526 => x"00", -- $0fc0e
          64527 => x"00", -- $0fc0f
          64528 => x"00", -- $0fc10
          64529 => x"00", -- $0fc11
          64530 => x"00", -- $0fc12
          64531 => x"00", -- $0fc13
          64532 => x"00", -- $0fc14
          64533 => x"00", -- $0fc15
          64534 => x"00", -- $0fc16
          64535 => x"00", -- $0fc17
          64536 => x"00", -- $0fc18
          64537 => x"00", -- $0fc19
          64538 => x"00", -- $0fc1a
          64539 => x"00", -- $0fc1b
          64540 => x"00", -- $0fc1c
          64541 => x"00", -- $0fc1d
          64542 => x"00", -- $0fc1e
          64543 => x"00", -- $0fc1f
          64544 => x"00", -- $0fc20
          64545 => x"00", -- $0fc21
          64546 => x"00", -- $0fc22
          64547 => x"00", -- $0fc23
          64548 => x"00", -- $0fc24
          64549 => x"00", -- $0fc25
          64550 => x"00", -- $0fc26
          64551 => x"00", -- $0fc27
          64552 => x"00", -- $0fc28
          64553 => x"00", -- $0fc29
          64554 => x"00", -- $0fc2a
          64555 => x"00", -- $0fc2b
          64556 => x"00", -- $0fc2c
          64557 => x"00", -- $0fc2d
          64558 => x"00", -- $0fc2e
          64559 => x"00", -- $0fc2f
          64560 => x"00", -- $0fc30
          64561 => x"00", -- $0fc31
          64562 => x"00", -- $0fc32
          64563 => x"00", -- $0fc33
          64564 => x"00", -- $0fc34
          64565 => x"00", -- $0fc35
          64566 => x"00", -- $0fc36
          64567 => x"00", -- $0fc37
          64568 => x"00", -- $0fc38
          64569 => x"00", -- $0fc39
          64570 => x"00", -- $0fc3a
          64571 => x"00", -- $0fc3b
          64572 => x"00", -- $0fc3c
          64573 => x"00", -- $0fc3d
          64574 => x"00", -- $0fc3e
          64575 => x"00", -- $0fc3f
          64576 => x"00", -- $0fc40
          64577 => x"00", -- $0fc41
          64578 => x"00", -- $0fc42
          64579 => x"00", -- $0fc43
          64580 => x"00", -- $0fc44
          64581 => x"00", -- $0fc45
          64582 => x"00", -- $0fc46
          64583 => x"00", -- $0fc47
          64584 => x"00", -- $0fc48
          64585 => x"00", -- $0fc49
          64586 => x"00", -- $0fc4a
          64587 => x"00", -- $0fc4b
          64588 => x"00", -- $0fc4c
          64589 => x"00", -- $0fc4d
          64590 => x"00", -- $0fc4e
          64591 => x"00", -- $0fc4f
          64592 => x"00", -- $0fc50
          64593 => x"00", -- $0fc51
          64594 => x"00", -- $0fc52
          64595 => x"00", -- $0fc53
          64596 => x"00", -- $0fc54
          64597 => x"00", -- $0fc55
          64598 => x"00", -- $0fc56
          64599 => x"00", -- $0fc57
          64600 => x"00", -- $0fc58
          64601 => x"00", -- $0fc59
          64602 => x"00", -- $0fc5a
          64603 => x"00", -- $0fc5b
          64604 => x"00", -- $0fc5c
          64605 => x"00", -- $0fc5d
          64606 => x"00", -- $0fc5e
          64607 => x"00", -- $0fc5f
          64608 => x"00", -- $0fc60
          64609 => x"00", -- $0fc61
          64610 => x"00", -- $0fc62
          64611 => x"00", -- $0fc63
          64612 => x"00", -- $0fc64
          64613 => x"00", -- $0fc65
          64614 => x"00", -- $0fc66
          64615 => x"00", -- $0fc67
          64616 => x"00", -- $0fc68
          64617 => x"00", -- $0fc69
          64618 => x"00", -- $0fc6a
          64619 => x"00", -- $0fc6b
          64620 => x"00", -- $0fc6c
          64621 => x"00", -- $0fc6d
          64622 => x"00", -- $0fc6e
          64623 => x"00", -- $0fc6f
          64624 => x"00", -- $0fc70
          64625 => x"00", -- $0fc71
          64626 => x"00", -- $0fc72
          64627 => x"00", -- $0fc73
          64628 => x"00", -- $0fc74
          64629 => x"00", -- $0fc75
          64630 => x"00", -- $0fc76
          64631 => x"00", -- $0fc77
          64632 => x"00", -- $0fc78
          64633 => x"00", -- $0fc79
          64634 => x"00", -- $0fc7a
          64635 => x"00", -- $0fc7b
          64636 => x"00", -- $0fc7c
          64637 => x"00", -- $0fc7d
          64638 => x"00", -- $0fc7e
          64639 => x"00", -- $0fc7f
          64640 => x"00", -- $0fc80
          64641 => x"00", -- $0fc81
          64642 => x"00", -- $0fc82
          64643 => x"00", -- $0fc83
          64644 => x"00", -- $0fc84
          64645 => x"00", -- $0fc85
          64646 => x"00", -- $0fc86
          64647 => x"00", -- $0fc87
          64648 => x"00", -- $0fc88
          64649 => x"00", -- $0fc89
          64650 => x"00", -- $0fc8a
          64651 => x"00", -- $0fc8b
          64652 => x"00", -- $0fc8c
          64653 => x"00", -- $0fc8d
          64654 => x"00", -- $0fc8e
          64655 => x"00", -- $0fc8f
          64656 => x"00", -- $0fc90
          64657 => x"00", -- $0fc91
          64658 => x"00", -- $0fc92
          64659 => x"00", -- $0fc93
          64660 => x"00", -- $0fc94
          64661 => x"00", -- $0fc95
          64662 => x"00", -- $0fc96
          64663 => x"00", -- $0fc97
          64664 => x"00", -- $0fc98
          64665 => x"00", -- $0fc99
          64666 => x"00", -- $0fc9a
          64667 => x"00", -- $0fc9b
          64668 => x"00", -- $0fc9c
          64669 => x"00", -- $0fc9d
          64670 => x"00", -- $0fc9e
          64671 => x"00", -- $0fc9f
          64672 => x"00", -- $0fca0
          64673 => x"00", -- $0fca1
          64674 => x"00", -- $0fca2
          64675 => x"00", -- $0fca3
          64676 => x"00", -- $0fca4
          64677 => x"00", -- $0fca5
          64678 => x"00", -- $0fca6
          64679 => x"00", -- $0fca7
          64680 => x"00", -- $0fca8
          64681 => x"00", -- $0fca9
          64682 => x"00", -- $0fcaa
          64683 => x"00", -- $0fcab
          64684 => x"00", -- $0fcac
          64685 => x"00", -- $0fcad
          64686 => x"00", -- $0fcae
          64687 => x"00", -- $0fcaf
          64688 => x"00", -- $0fcb0
          64689 => x"00", -- $0fcb1
          64690 => x"00", -- $0fcb2
          64691 => x"00", -- $0fcb3
          64692 => x"00", -- $0fcb4
          64693 => x"00", -- $0fcb5
          64694 => x"00", -- $0fcb6
          64695 => x"00", -- $0fcb7
          64696 => x"00", -- $0fcb8
          64697 => x"00", -- $0fcb9
          64698 => x"00", -- $0fcba
          64699 => x"00", -- $0fcbb
          64700 => x"00", -- $0fcbc
          64701 => x"00", -- $0fcbd
          64702 => x"00", -- $0fcbe
          64703 => x"00", -- $0fcbf
          64704 => x"00", -- $0fcc0
          64705 => x"00", -- $0fcc1
          64706 => x"00", -- $0fcc2
          64707 => x"00", -- $0fcc3
          64708 => x"00", -- $0fcc4
          64709 => x"00", -- $0fcc5
          64710 => x"00", -- $0fcc6
          64711 => x"00", -- $0fcc7
          64712 => x"00", -- $0fcc8
          64713 => x"00", -- $0fcc9
          64714 => x"00", -- $0fcca
          64715 => x"00", -- $0fccb
          64716 => x"00", -- $0fccc
          64717 => x"00", -- $0fccd
          64718 => x"00", -- $0fcce
          64719 => x"00", -- $0fccf
          64720 => x"00", -- $0fcd0
          64721 => x"00", -- $0fcd1
          64722 => x"00", -- $0fcd2
          64723 => x"00", -- $0fcd3
          64724 => x"00", -- $0fcd4
          64725 => x"00", -- $0fcd5
          64726 => x"00", -- $0fcd6
          64727 => x"00", -- $0fcd7
          64728 => x"00", -- $0fcd8
          64729 => x"00", -- $0fcd9
          64730 => x"00", -- $0fcda
          64731 => x"00", -- $0fcdb
          64732 => x"00", -- $0fcdc
          64733 => x"00", -- $0fcdd
          64734 => x"00", -- $0fcde
          64735 => x"00", -- $0fcdf
          64736 => x"00", -- $0fce0
          64737 => x"00", -- $0fce1
          64738 => x"00", -- $0fce2
          64739 => x"00", -- $0fce3
          64740 => x"00", -- $0fce4
          64741 => x"00", -- $0fce5
          64742 => x"00", -- $0fce6
          64743 => x"00", -- $0fce7
          64744 => x"00", -- $0fce8
          64745 => x"00", -- $0fce9
          64746 => x"00", -- $0fcea
          64747 => x"00", -- $0fceb
          64748 => x"00", -- $0fcec
          64749 => x"00", -- $0fced
          64750 => x"00", -- $0fcee
          64751 => x"00", -- $0fcef
          64752 => x"00", -- $0fcf0
          64753 => x"00", -- $0fcf1
          64754 => x"00", -- $0fcf2
          64755 => x"00", -- $0fcf3
          64756 => x"00", -- $0fcf4
          64757 => x"00", -- $0fcf5
          64758 => x"00", -- $0fcf6
          64759 => x"00", -- $0fcf7
          64760 => x"00", -- $0fcf8
          64761 => x"00", -- $0fcf9
          64762 => x"00", -- $0fcfa
          64763 => x"00", -- $0fcfb
          64764 => x"00", -- $0fcfc
          64765 => x"00", -- $0fcfd
          64766 => x"00", -- $0fcfe
          64767 => x"00", -- $0fcff
          64768 => x"00", -- $0fd00
          64769 => x"00", -- $0fd01
          64770 => x"00", -- $0fd02
          64771 => x"00", -- $0fd03
          64772 => x"00", -- $0fd04
          64773 => x"00", -- $0fd05
          64774 => x"00", -- $0fd06
          64775 => x"00", -- $0fd07
          64776 => x"00", -- $0fd08
          64777 => x"00", -- $0fd09
          64778 => x"00", -- $0fd0a
          64779 => x"00", -- $0fd0b
          64780 => x"00", -- $0fd0c
          64781 => x"00", -- $0fd0d
          64782 => x"00", -- $0fd0e
          64783 => x"00", -- $0fd0f
          64784 => x"00", -- $0fd10
          64785 => x"00", -- $0fd11
          64786 => x"00", -- $0fd12
          64787 => x"00", -- $0fd13
          64788 => x"00", -- $0fd14
          64789 => x"00", -- $0fd15
          64790 => x"00", -- $0fd16
          64791 => x"00", -- $0fd17
          64792 => x"00", -- $0fd18
          64793 => x"00", -- $0fd19
          64794 => x"00", -- $0fd1a
          64795 => x"00", -- $0fd1b
          64796 => x"00", -- $0fd1c
          64797 => x"00", -- $0fd1d
          64798 => x"00", -- $0fd1e
          64799 => x"00", -- $0fd1f
          64800 => x"00", -- $0fd20
          64801 => x"00", -- $0fd21
          64802 => x"00", -- $0fd22
          64803 => x"00", -- $0fd23
          64804 => x"00", -- $0fd24
          64805 => x"00", -- $0fd25
          64806 => x"00", -- $0fd26
          64807 => x"00", -- $0fd27
          64808 => x"00", -- $0fd28
          64809 => x"00", -- $0fd29
          64810 => x"00", -- $0fd2a
          64811 => x"00", -- $0fd2b
          64812 => x"00", -- $0fd2c
          64813 => x"00", -- $0fd2d
          64814 => x"00", -- $0fd2e
          64815 => x"00", -- $0fd2f
          64816 => x"00", -- $0fd30
          64817 => x"00", -- $0fd31
          64818 => x"00", -- $0fd32
          64819 => x"00", -- $0fd33
          64820 => x"00", -- $0fd34
          64821 => x"00", -- $0fd35
          64822 => x"00", -- $0fd36
          64823 => x"00", -- $0fd37
          64824 => x"00", -- $0fd38
          64825 => x"00", -- $0fd39
          64826 => x"00", -- $0fd3a
          64827 => x"00", -- $0fd3b
          64828 => x"00", -- $0fd3c
          64829 => x"00", -- $0fd3d
          64830 => x"00", -- $0fd3e
          64831 => x"00", -- $0fd3f
          64832 => x"00", -- $0fd40
          64833 => x"00", -- $0fd41
          64834 => x"00", -- $0fd42
          64835 => x"00", -- $0fd43
          64836 => x"00", -- $0fd44
          64837 => x"00", -- $0fd45
          64838 => x"00", -- $0fd46
          64839 => x"00", -- $0fd47
          64840 => x"00", -- $0fd48
          64841 => x"00", -- $0fd49
          64842 => x"00", -- $0fd4a
          64843 => x"00", -- $0fd4b
          64844 => x"00", -- $0fd4c
          64845 => x"00", -- $0fd4d
          64846 => x"00", -- $0fd4e
          64847 => x"00", -- $0fd4f
          64848 => x"00", -- $0fd50
          64849 => x"00", -- $0fd51
          64850 => x"00", -- $0fd52
          64851 => x"00", -- $0fd53
          64852 => x"00", -- $0fd54
          64853 => x"00", -- $0fd55
          64854 => x"00", -- $0fd56
          64855 => x"00", -- $0fd57
          64856 => x"00", -- $0fd58
          64857 => x"00", -- $0fd59
          64858 => x"00", -- $0fd5a
          64859 => x"00", -- $0fd5b
          64860 => x"00", -- $0fd5c
          64861 => x"00", -- $0fd5d
          64862 => x"00", -- $0fd5e
          64863 => x"00", -- $0fd5f
          64864 => x"00", -- $0fd60
          64865 => x"00", -- $0fd61
          64866 => x"00", -- $0fd62
          64867 => x"00", -- $0fd63
          64868 => x"00", -- $0fd64
          64869 => x"00", -- $0fd65
          64870 => x"00", -- $0fd66
          64871 => x"00", -- $0fd67
          64872 => x"00", -- $0fd68
          64873 => x"00", -- $0fd69
          64874 => x"00", -- $0fd6a
          64875 => x"00", -- $0fd6b
          64876 => x"00", -- $0fd6c
          64877 => x"00", -- $0fd6d
          64878 => x"00", -- $0fd6e
          64879 => x"00", -- $0fd6f
          64880 => x"00", -- $0fd70
          64881 => x"00", -- $0fd71
          64882 => x"00", -- $0fd72
          64883 => x"00", -- $0fd73
          64884 => x"00", -- $0fd74
          64885 => x"00", -- $0fd75
          64886 => x"00", -- $0fd76
          64887 => x"00", -- $0fd77
          64888 => x"00", -- $0fd78
          64889 => x"00", -- $0fd79
          64890 => x"00", -- $0fd7a
          64891 => x"00", -- $0fd7b
          64892 => x"00", -- $0fd7c
          64893 => x"00", -- $0fd7d
          64894 => x"00", -- $0fd7e
          64895 => x"00", -- $0fd7f
          64896 => x"00", -- $0fd80
          64897 => x"00", -- $0fd81
          64898 => x"00", -- $0fd82
          64899 => x"00", -- $0fd83
          64900 => x"00", -- $0fd84
          64901 => x"00", -- $0fd85
          64902 => x"00", -- $0fd86
          64903 => x"00", -- $0fd87
          64904 => x"00", -- $0fd88
          64905 => x"00", -- $0fd89
          64906 => x"00", -- $0fd8a
          64907 => x"00", -- $0fd8b
          64908 => x"00", -- $0fd8c
          64909 => x"00", -- $0fd8d
          64910 => x"00", -- $0fd8e
          64911 => x"00", -- $0fd8f
          64912 => x"00", -- $0fd90
          64913 => x"00", -- $0fd91
          64914 => x"00", -- $0fd92
          64915 => x"00", -- $0fd93
          64916 => x"00", -- $0fd94
          64917 => x"00", -- $0fd95
          64918 => x"00", -- $0fd96
          64919 => x"00", -- $0fd97
          64920 => x"00", -- $0fd98
          64921 => x"00", -- $0fd99
          64922 => x"00", -- $0fd9a
          64923 => x"00", -- $0fd9b
          64924 => x"00", -- $0fd9c
          64925 => x"00", -- $0fd9d
          64926 => x"00", -- $0fd9e
          64927 => x"00", -- $0fd9f
          64928 => x"00", -- $0fda0
          64929 => x"00", -- $0fda1
          64930 => x"00", -- $0fda2
          64931 => x"00", -- $0fda3
          64932 => x"00", -- $0fda4
          64933 => x"00", -- $0fda5
          64934 => x"00", -- $0fda6
          64935 => x"00", -- $0fda7
          64936 => x"00", -- $0fda8
          64937 => x"00", -- $0fda9
          64938 => x"00", -- $0fdaa
          64939 => x"00", -- $0fdab
          64940 => x"00", -- $0fdac
          64941 => x"00", -- $0fdad
          64942 => x"00", -- $0fdae
          64943 => x"00", -- $0fdaf
          64944 => x"00", -- $0fdb0
          64945 => x"00", -- $0fdb1
          64946 => x"00", -- $0fdb2
          64947 => x"00", -- $0fdb3
          64948 => x"00", -- $0fdb4
          64949 => x"00", -- $0fdb5
          64950 => x"00", -- $0fdb6
          64951 => x"00", -- $0fdb7
          64952 => x"00", -- $0fdb8
          64953 => x"00", -- $0fdb9
          64954 => x"00", -- $0fdba
          64955 => x"00", -- $0fdbb
          64956 => x"00", -- $0fdbc
          64957 => x"00", -- $0fdbd
          64958 => x"00", -- $0fdbe
          64959 => x"00", -- $0fdbf
          64960 => x"00", -- $0fdc0
          64961 => x"00", -- $0fdc1
          64962 => x"00", -- $0fdc2
          64963 => x"00", -- $0fdc3
          64964 => x"00", -- $0fdc4
          64965 => x"00", -- $0fdc5
          64966 => x"00", -- $0fdc6
          64967 => x"00", -- $0fdc7
          64968 => x"00", -- $0fdc8
          64969 => x"00", -- $0fdc9
          64970 => x"00", -- $0fdca
          64971 => x"00", -- $0fdcb
          64972 => x"00", -- $0fdcc
          64973 => x"00", -- $0fdcd
          64974 => x"00", -- $0fdce
          64975 => x"00", -- $0fdcf
          64976 => x"00", -- $0fdd0
          64977 => x"00", -- $0fdd1
          64978 => x"00", -- $0fdd2
          64979 => x"00", -- $0fdd3
          64980 => x"00", -- $0fdd4
          64981 => x"00", -- $0fdd5
          64982 => x"00", -- $0fdd6
          64983 => x"00", -- $0fdd7
          64984 => x"00", -- $0fdd8
          64985 => x"00", -- $0fdd9
          64986 => x"00", -- $0fdda
          64987 => x"00", -- $0fddb
          64988 => x"00", -- $0fddc
          64989 => x"00", -- $0fddd
          64990 => x"00", -- $0fdde
          64991 => x"00", -- $0fddf
          64992 => x"00", -- $0fde0
          64993 => x"00", -- $0fde1
          64994 => x"00", -- $0fde2
          64995 => x"00", -- $0fde3
          64996 => x"00", -- $0fde4
          64997 => x"00", -- $0fde5
          64998 => x"00", -- $0fde6
          64999 => x"00", -- $0fde7
          65000 => x"00", -- $0fde8
          65001 => x"00", -- $0fde9
          65002 => x"00", -- $0fdea
          65003 => x"00", -- $0fdeb
          65004 => x"00", -- $0fdec
          65005 => x"00", -- $0fded
          65006 => x"00", -- $0fdee
          65007 => x"00", -- $0fdef
          65008 => x"00", -- $0fdf0
          65009 => x"00", -- $0fdf1
          65010 => x"00", -- $0fdf2
          65011 => x"00", -- $0fdf3
          65012 => x"00", -- $0fdf4
          65013 => x"00", -- $0fdf5
          65014 => x"00", -- $0fdf6
          65015 => x"00", -- $0fdf7
          65016 => x"00", -- $0fdf8
          65017 => x"00", -- $0fdf9
          65018 => x"00", -- $0fdfa
          65019 => x"00", -- $0fdfb
          65020 => x"00", -- $0fdfc
          65021 => x"00", -- $0fdfd
          65022 => x"00", -- $0fdfe
          65023 => x"00", -- $0fdff
          65024 => x"00", -- $0fe00
          65025 => x"00", -- $0fe01
          65026 => x"00", -- $0fe02
          65027 => x"00", -- $0fe03
          65028 => x"00", -- $0fe04
          65029 => x"00", -- $0fe05
          65030 => x"00", -- $0fe06
          65031 => x"00", -- $0fe07
          65032 => x"00", -- $0fe08
          65033 => x"00", -- $0fe09
          65034 => x"00", -- $0fe0a
          65035 => x"00", -- $0fe0b
          65036 => x"00", -- $0fe0c
          65037 => x"00", -- $0fe0d
          65038 => x"00", -- $0fe0e
          65039 => x"00", -- $0fe0f
          65040 => x"00", -- $0fe10
          65041 => x"00", -- $0fe11
          65042 => x"00", -- $0fe12
          65043 => x"00", -- $0fe13
          65044 => x"00", -- $0fe14
          65045 => x"00", -- $0fe15
          65046 => x"00", -- $0fe16
          65047 => x"00", -- $0fe17
          65048 => x"00", -- $0fe18
          65049 => x"00", -- $0fe19
          65050 => x"00", -- $0fe1a
          65051 => x"00", -- $0fe1b
          65052 => x"00", -- $0fe1c
          65053 => x"00", -- $0fe1d
          65054 => x"00", -- $0fe1e
          65055 => x"00", -- $0fe1f
          65056 => x"00", -- $0fe20
          65057 => x"00", -- $0fe21
          65058 => x"00", -- $0fe22
          65059 => x"00", -- $0fe23
          65060 => x"00", -- $0fe24
          65061 => x"00", -- $0fe25
          65062 => x"00", -- $0fe26
          65063 => x"00", -- $0fe27
          65064 => x"00", -- $0fe28
          65065 => x"00", -- $0fe29
          65066 => x"00", -- $0fe2a
          65067 => x"00", -- $0fe2b
          65068 => x"00", -- $0fe2c
          65069 => x"00", -- $0fe2d
          65070 => x"00", -- $0fe2e
          65071 => x"00", -- $0fe2f
          65072 => x"00", -- $0fe30
          65073 => x"00", -- $0fe31
          65074 => x"00", -- $0fe32
          65075 => x"00", -- $0fe33
          65076 => x"00", -- $0fe34
          65077 => x"00", -- $0fe35
          65078 => x"00", -- $0fe36
          65079 => x"00", -- $0fe37
          65080 => x"00", -- $0fe38
          65081 => x"00", -- $0fe39
          65082 => x"00", -- $0fe3a
          65083 => x"00", -- $0fe3b
          65084 => x"00", -- $0fe3c
          65085 => x"00", -- $0fe3d
          65086 => x"00", -- $0fe3e
          65087 => x"00", -- $0fe3f
          65088 => x"00", -- $0fe40
          65089 => x"00", -- $0fe41
          65090 => x"00", -- $0fe42
          65091 => x"00", -- $0fe43
          65092 => x"00", -- $0fe44
          65093 => x"00", -- $0fe45
          65094 => x"00", -- $0fe46
          65095 => x"00", -- $0fe47
          65096 => x"00", -- $0fe48
          65097 => x"00", -- $0fe49
          65098 => x"00", -- $0fe4a
          65099 => x"00", -- $0fe4b
          65100 => x"00", -- $0fe4c
          65101 => x"00", -- $0fe4d
          65102 => x"00", -- $0fe4e
          65103 => x"00", -- $0fe4f
          65104 => x"00", -- $0fe50
          65105 => x"00", -- $0fe51
          65106 => x"00", -- $0fe52
          65107 => x"00", -- $0fe53
          65108 => x"00", -- $0fe54
          65109 => x"00", -- $0fe55
          65110 => x"00", -- $0fe56
          65111 => x"00", -- $0fe57
          65112 => x"00", -- $0fe58
          65113 => x"00", -- $0fe59
          65114 => x"00", -- $0fe5a
          65115 => x"00", -- $0fe5b
          65116 => x"00", -- $0fe5c
          65117 => x"00", -- $0fe5d
          65118 => x"00", -- $0fe5e
          65119 => x"00", -- $0fe5f
          65120 => x"00", -- $0fe60
          65121 => x"00", -- $0fe61
          65122 => x"00", -- $0fe62
          65123 => x"00", -- $0fe63
          65124 => x"00", -- $0fe64
          65125 => x"00", -- $0fe65
          65126 => x"00", -- $0fe66
          65127 => x"00", -- $0fe67
          65128 => x"00", -- $0fe68
          65129 => x"00", -- $0fe69
          65130 => x"00", -- $0fe6a
          65131 => x"00", -- $0fe6b
          65132 => x"00", -- $0fe6c
          65133 => x"00", -- $0fe6d
          65134 => x"00", -- $0fe6e
          65135 => x"00", -- $0fe6f
          65136 => x"00", -- $0fe70
          65137 => x"00", -- $0fe71
          65138 => x"00", -- $0fe72
          65139 => x"00", -- $0fe73
          65140 => x"00", -- $0fe74
          65141 => x"00", -- $0fe75
          65142 => x"00", -- $0fe76
          65143 => x"00", -- $0fe77
          65144 => x"00", -- $0fe78
          65145 => x"00", -- $0fe79
          65146 => x"00", -- $0fe7a
          65147 => x"00", -- $0fe7b
          65148 => x"00", -- $0fe7c
          65149 => x"00", -- $0fe7d
          65150 => x"00", -- $0fe7e
          65151 => x"00", -- $0fe7f
          65152 => x"00", -- $0fe80
          65153 => x"00", -- $0fe81
          65154 => x"00", -- $0fe82
          65155 => x"00", -- $0fe83
          65156 => x"00", -- $0fe84
          65157 => x"00", -- $0fe85
          65158 => x"00", -- $0fe86
          65159 => x"00", -- $0fe87
          65160 => x"00", -- $0fe88
          65161 => x"00", -- $0fe89
          65162 => x"00", -- $0fe8a
          65163 => x"00", -- $0fe8b
          65164 => x"00", -- $0fe8c
          65165 => x"00", -- $0fe8d
          65166 => x"00", -- $0fe8e
          65167 => x"00", -- $0fe8f
          65168 => x"00", -- $0fe90
          65169 => x"00", -- $0fe91
          65170 => x"00", -- $0fe92
          65171 => x"00", -- $0fe93
          65172 => x"00", -- $0fe94
          65173 => x"00", -- $0fe95
          65174 => x"00", -- $0fe96
          65175 => x"00", -- $0fe97
          65176 => x"00", -- $0fe98
          65177 => x"00", -- $0fe99
          65178 => x"00", -- $0fe9a
          65179 => x"00", -- $0fe9b
          65180 => x"00", -- $0fe9c
          65181 => x"00", -- $0fe9d
          65182 => x"00", -- $0fe9e
          65183 => x"00", -- $0fe9f
          65184 => x"00", -- $0fea0
          65185 => x"00", -- $0fea1
          65186 => x"00", -- $0fea2
          65187 => x"00", -- $0fea3
          65188 => x"00", -- $0fea4
          65189 => x"00", -- $0fea5
          65190 => x"00", -- $0fea6
          65191 => x"00", -- $0fea7
          65192 => x"00", -- $0fea8
          65193 => x"00", -- $0fea9
          65194 => x"00", -- $0feaa
          65195 => x"00", -- $0feab
          65196 => x"00", -- $0feac
          65197 => x"00", -- $0fead
          65198 => x"00", -- $0feae
          65199 => x"00", -- $0feaf
          65200 => x"00", -- $0feb0
          65201 => x"00", -- $0feb1
          65202 => x"00", -- $0feb2
          65203 => x"00", -- $0feb3
          65204 => x"00", -- $0feb4
          65205 => x"00", -- $0feb5
          65206 => x"00", -- $0feb6
          65207 => x"00", -- $0feb7
          65208 => x"00", -- $0feb8
          65209 => x"00", -- $0feb9
          65210 => x"00", -- $0feba
          65211 => x"00", -- $0febb
          65212 => x"00", -- $0febc
          65213 => x"00", -- $0febd
          65214 => x"00", -- $0febe
          65215 => x"00", -- $0febf
          65216 => x"00", -- $0fec0
          65217 => x"00", -- $0fec1
          65218 => x"00", -- $0fec2
          65219 => x"00", -- $0fec3
          65220 => x"00", -- $0fec4
          65221 => x"00", -- $0fec5
          65222 => x"00", -- $0fec6
          65223 => x"00", -- $0fec7
          65224 => x"00", -- $0fec8
          65225 => x"00", -- $0fec9
          65226 => x"00", -- $0feca
          65227 => x"00", -- $0fecb
          65228 => x"00", -- $0fecc
          65229 => x"00", -- $0fecd
          65230 => x"00", -- $0fece
          65231 => x"00", -- $0fecf
          65232 => x"00", -- $0fed0
          65233 => x"00", -- $0fed1
          65234 => x"00", -- $0fed2
          65235 => x"00", -- $0fed3
          65236 => x"00", -- $0fed4
          65237 => x"00", -- $0fed5
          65238 => x"00", -- $0fed6
          65239 => x"00", -- $0fed7
          65240 => x"00", -- $0fed8
          65241 => x"00", -- $0fed9
          65242 => x"00", -- $0feda
          65243 => x"00", -- $0fedb
          65244 => x"00", -- $0fedc
          65245 => x"00", -- $0fedd
          65246 => x"00", -- $0fede
          65247 => x"00", -- $0fedf
          65248 => x"00", -- $0fee0
          65249 => x"00", -- $0fee1
          65250 => x"00", -- $0fee2
          65251 => x"00", -- $0fee3
          65252 => x"00", -- $0fee4
          65253 => x"00", -- $0fee5
          65254 => x"00", -- $0fee6
          65255 => x"00", -- $0fee7
          65256 => x"00", -- $0fee8
          65257 => x"00", -- $0fee9
          65258 => x"00", -- $0feea
          65259 => x"00", -- $0feeb
          65260 => x"00", -- $0feec
          65261 => x"00", -- $0feed
          65262 => x"00", -- $0feee
          65263 => x"00", -- $0feef
          65264 => x"00", -- $0fef0
          65265 => x"00", -- $0fef1
          65266 => x"00", -- $0fef2
          65267 => x"00", -- $0fef3
          65268 => x"00", -- $0fef4
          65269 => x"00", -- $0fef5
          65270 => x"00", -- $0fef6
          65271 => x"00", -- $0fef7
          65272 => x"00", -- $0fef8
          65273 => x"00", -- $0fef9
          65274 => x"00", -- $0fefa
          65275 => x"00", -- $0fefb
          65276 => x"00", -- $0fefc
          65277 => x"00", -- $0fefd
          65278 => x"00", -- $0fefe
          65279 => x"00", -- $0feff
          65280 => x"00", -- $0ff00
          65281 => x"00", -- $0ff01
          65282 => x"00", -- $0ff02
          65283 => x"00", -- $0ff03
          65284 => x"00", -- $0ff04
          65285 => x"00", -- $0ff05
          65286 => x"00", -- $0ff06
          65287 => x"00", -- $0ff07
          65288 => x"00", -- $0ff08
          65289 => x"00", -- $0ff09
          65290 => x"00", -- $0ff0a
          65291 => x"00", -- $0ff0b
          65292 => x"00", -- $0ff0c
          65293 => x"00", -- $0ff0d
          65294 => x"00", -- $0ff0e
          65295 => x"00", -- $0ff0f
          65296 => x"00", -- $0ff10
          65297 => x"00", -- $0ff11
          65298 => x"00", -- $0ff12
          65299 => x"00", -- $0ff13
          65300 => x"00", -- $0ff14
          65301 => x"00", -- $0ff15
          65302 => x"00", -- $0ff16
          65303 => x"00", -- $0ff17
          65304 => x"00", -- $0ff18
          65305 => x"00", -- $0ff19
          65306 => x"00", -- $0ff1a
          65307 => x"00", -- $0ff1b
          65308 => x"00", -- $0ff1c
          65309 => x"00", -- $0ff1d
          65310 => x"00", -- $0ff1e
          65311 => x"00", -- $0ff1f
          65312 => x"00", -- $0ff20
          65313 => x"00", -- $0ff21
          65314 => x"00", -- $0ff22
          65315 => x"00", -- $0ff23
          65316 => x"00", -- $0ff24
          65317 => x"00", -- $0ff25
          65318 => x"00", -- $0ff26
          65319 => x"00", -- $0ff27
          65320 => x"00", -- $0ff28
          65321 => x"00", -- $0ff29
          65322 => x"00", -- $0ff2a
          65323 => x"00", -- $0ff2b
          65324 => x"00", -- $0ff2c
          65325 => x"00", -- $0ff2d
          65326 => x"00", -- $0ff2e
          65327 => x"00", -- $0ff2f
          65328 => x"00", -- $0ff30
          65329 => x"00", -- $0ff31
          65330 => x"00", -- $0ff32
          65331 => x"00", -- $0ff33
          65332 => x"00", -- $0ff34
          65333 => x"00", -- $0ff35
          65334 => x"00", -- $0ff36
          65335 => x"00", -- $0ff37
          65336 => x"00", -- $0ff38
          65337 => x"00", -- $0ff39
          65338 => x"00", -- $0ff3a
          65339 => x"00", -- $0ff3b
          65340 => x"00", -- $0ff3c
          65341 => x"00", -- $0ff3d
          65342 => x"00", -- $0ff3e
          65343 => x"00", -- $0ff3f
          65344 => x"00", -- $0ff40
          65345 => x"00", -- $0ff41
          65346 => x"00", -- $0ff42
          65347 => x"00", -- $0ff43
          65348 => x"00", -- $0ff44
          65349 => x"00", -- $0ff45
          65350 => x"00", -- $0ff46
          65351 => x"00", -- $0ff47
          65352 => x"00", -- $0ff48
          65353 => x"00", -- $0ff49
          65354 => x"00", -- $0ff4a
          65355 => x"00", -- $0ff4b
          65356 => x"00", -- $0ff4c
          65357 => x"00", -- $0ff4d
          65358 => x"00", -- $0ff4e
          65359 => x"00", -- $0ff4f
          65360 => x"00", -- $0ff50
          65361 => x"00", -- $0ff51
          65362 => x"00", -- $0ff52
          65363 => x"00", -- $0ff53
          65364 => x"00", -- $0ff54
          65365 => x"00", -- $0ff55
          65366 => x"00", -- $0ff56
          65367 => x"00", -- $0ff57
          65368 => x"00", -- $0ff58
          65369 => x"00", -- $0ff59
          65370 => x"00", -- $0ff5a
          65371 => x"00", -- $0ff5b
          65372 => x"00", -- $0ff5c
          65373 => x"00", -- $0ff5d
          65374 => x"00", -- $0ff5e
          65375 => x"00", -- $0ff5f
          65376 => x"00", -- $0ff60
          65377 => x"00", -- $0ff61
          65378 => x"00", -- $0ff62
          65379 => x"00", -- $0ff63
          65380 => x"00", -- $0ff64
          65381 => x"00", -- $0ff65
          65382 => x"00", -- $0ff66
          65383 => x"00", -- $0ff67
          65384 => x"00", -- $0ff68
          65385 => x"00", -- $0ff69
          65386 => x"00", -- $0ff6a
          65387 => x"00", -- $0ff6b
          65388 => x"00", -- $0ff6c
          65389 => x"00", -- $0ff6d
          65390 => x"00", -- $0ff6e
          65391 => x"00", -- $0ff6f
          65392 => x"00", -- $0ff70
          65393 => x"00", -- $0ff71
          65394 => x"00", -- $0ff72
          65395 => x"00", -- $0ff73
          65396 => x"00", -- $0ff74
          65397 => x"00", -- $0ff75
          65398 => x"00", -- $0ff76
          65399 => x"00", -- $0ff77
          65400 => x"00", -- $0ff78
          65401 => x"00", -- $0ff79
          65402 => x"00", -- $0ff7a
          65403 => x"00", -- $0ff7b
          65404 => x"00", -- $0ff7c
          65405 => x"00", -- $0ff7d
          65406 => x"00", -- $0ff7e
          65407 => x"00", -- $0ff7f
          65408 => x"00", -- $0ff80
          65409 => x"00", -- $0ff81
          65410 => x"00", -- $0ff82
          65411 => x"00", -- $0ff83
          65412 => x"00", -- $0ff84
          65413 => x"00", -- $0ff85
          65414 => x"00", -- $0ff86
          65415 => x"00", -- $0ff87
          65416 => x"00", -- $0ff88
          65417 => x"00", -- $0ff89
          65418 => x"00", -- $0ff8a
          65419 => x"00", -- $0ff8b
          65420 => x"00", -- $0ff8c
          65421 => x"00", -- $0ff8d
          65422 => x"00", -- $0ff8e
          65423 => x"00", -- $0ff8f
          65424 => x"00", -- $0ff90
          65425 => x"00", -- $0ff91
          65426 => x"00", -- $0ff92
          65427 => x"00", -- $0ff93
          65428 => x"00", -- $0ff94
          65429 => x"00", -- $0ff95
          65430 => x"00", -- $0ff96
          65431 => x"00", -- $0ff97
          65432 => x"00", -- $0ff98
          65433 => x"00", -- $0ff99
          65434 => x"00", -- $0ff9a
          65435 => x"00", -- $0ff9b
          65436 => x"00", -- $0ff9c
          65437 => x"00", -- $0ff9d
          65438 => x"00", -- $0ff9e
          65439 => x"00", -- $0ff9f
          65440 => x"00", -- $0ffa0
          65441 => x"00", -- $0ffa1
          65442 => x"00", -- $0ffa2
          65443 => x"00", -- $0ffa3
          65444 => x"00", -- $0ffa4
          65445 => x"00", -- $0ffa5
          65446 => x"00", -- $0ffa6
          65447 => x"00", -- $0ffa7
          65448 => x"00", -- $0ffa8
          65449 => x"00", -- $0ffa9
          65450 => x"00", -- $0ffaa
          65451 => x"00", -- $0ffab
          65452 => x"00", -- $0ffac
          65453 => x"00", -- $0ffad
          65454 => x"00", -- $0ffae
          65455 => x"00", -- $0ffaf
          65456 => x"00", -- $0ffb0
          65457 => x"00", -- $0ffb1
          65458 => x"00", -- $0ffb2
          65459 => x"00", -- $0ffb3
          65460 => x"00", -- $0ffb4
          65461 => x"00", -- $0ffb5
          65462 => x"00", -- $0ffb6
          65463 => x"00", -- $0ffb7
          65464 => x"00", -- $0ffb8
          65465 => x"00", -- $0ffb9
          65466 => x"00", -- $0ffba
          65467 => x"00", -- $0ffbb
          65468 => x"00", -- $0ffbc
          65469 => x"00", -- $0ffbd
          65470 => x"00", -- $0ffbe
          65471 => x"00", -- $0ffbf
          65472 => x"00", -- $0ffc0
          65473 => x"00", -- $0ffc1
          65474 => x"00", -- $0ffc2
          65475 => x"00", -- $0ffc3
          65476 => x"00", -- $0ffc4
          65477 => x"00", -- $0ffc5
          65478 => x"00", -- $0ffc6
          65479 => x"00", -- $0ffc7
          65480 => x"00", -- $0ffc8
          65481 => x"00", -- $0ffc9
          65482 => x"00", -- $0ffca
          65483 => x"00", -- $0ffcb
          65484 => x"00", -- $0ffcc
          65485 => x"00", -- $0ffcd
          65486 => x"00", -- $0ffce
          65487 => x"00", -- $0ffcf
          65488 => x"00", -- $0ffd0
          65489 => x"00", -- $0ffd1
          65490 => x"00", -- $0ffd2
          65491 => x"00", -- $0ffd3
          65492 => x"00", -- $0ffd4
          65493 => x"00", -- $0ffd5
          65494 => x"00", -- $0ffd6
          65495 => x"00", -- $0ffd7
          65496 => x"00", -- $0ffd8
          65497 => x"00", -- $0ffd9
          65498 => x"00", -- $0ffda
          65499 => x"00", -- $0ffdb
          65500 => x"00", -- $0ffdc
          65501 => x"00", -- $0ffdd
          65502 => x"00", -- $0ffde
          65503 => x"00", -- $0ffdf
          65504 => x"00", -- $0ffe0
          65505 => x"00", -- $0ffe1
          65506 => x"00", -- $0ffe2
          65507 => x"00", -- $0ffe3
          65508 => x"00", -- $0ffe4
          65509 => x"00", -- $0ffe5
          65510 => x"00", -- $0ffe6
          65511 => x"00", -- $0ffe7
          65512 => x"00", -- $0ffe8
          65513 => x"00", -- $0ffe9
          65514 => x"00", -- $0ffea
          65515 => x"00", -- $0ffeb
          65516 => x"00", -- $0ffec
          65517 => x"00", -- $0ffed
          65518 => x"00", -- $0ffee
          65519 => x"00", -- $0ffef
          65520 => x"00", -- $0fff0
          65521 => x"00", -- $0fff1
          65522 => x"00", -- $0fff2
          65523 => x"00", -- $0fff3
          65524 => x"00", -- $0fff4
          65525 => x"00", -- $0fff5
          65526 => x"00", -- $0fff6
          65527 => x"00", -- $0fff7
          65528 => x"00", -- $0fff8
          65529 => x"00", -- $0fff9
          65530 => x"00", -- $0fffa
          65531 => x"00", -- $0fffb
          65532 => x"00", -- $0fffc
          65533 => x"00", -- $0fffd
          65534 => x"00", -- $0fffe
          65535 => x"00" -- $0ffff
          ); -- $10000
begin

--process for read and write operation.
  PROCESS(ClkA)
  BEGIN
    if(rising_edge(ClkA)) then 
        doa <= ram(addressa);
    end if;
  END PROCESS;

end Behavioral;
